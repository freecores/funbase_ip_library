--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity a2h_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal a2h_avalon_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal a2h_avalon_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal a2h_avalon_slave_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal a2h_avalon_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal a2h_avalon_slave_read : OUT STD_LOGIC;
                 signal a2h_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal a2h_avalon_slave_reset_n : OUT STD_LOGIC;
                 signal a2h_avalon_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal a2h_avalon_slave_write : OUT STD_LOGIC;
                 signal a2h_avalon_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_a2h_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave : OUT STD_LOGIC
              );
end entity a2h_avalon_slave_arbitrator;


architecture europa of a2h_avalon_slave_arbitrator is
                signal a2h_avalon_slave_allgrants :  STD_LOGIC;
                signal a2h_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal a2h_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal a2h_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal a2h_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal a2h_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal a2h_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal a2h_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal a2h_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal a2h_avalon_slave_begins_xfer :  STD_LOGIC;
                signal a2h_avalon_slave_end_xfer :  STD_LOGIC;
                signal a2h_avalon_slave_firsttransfer :  STD_LOGIC;
                signal a2h_avalon_slave_grant_vector :  STD_LOGIC;
                signal a2h_avalon_slave_in_a_read_cycle :  STD_LOGIC;
                signal a2h_avalon_slave_in_a_write_cycle :  STD_LOGIC;
                signal a2h_avalon_slave_master_qreq_vector :  STD_LOGIC;
                signal a2h_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal a2h_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal a2h_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal a2h_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal a2h_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal a2h_avalon_slave_waits_for_read :  STD_LOGIC;
                signal a2h_avalon_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_a2h_avalon_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_a2h_avalon_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_saved_grant_a2h_avalon_slave :  STD_LOGIC;
                signal shifted_address_to_a2h_avalon_slave_from_pcie_to_hibi_4x_sopc_burst_5_downstream :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_a2h_avalon_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT a2h_avalon_slave_end_xfer;
    end if;

  end process;

  a2h_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave);
  --assign a2h_avalon_slave_readdata_from_sa = a2h_avalon_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  a2h_avalon_slave_readdata_from_sa <= a2h_avalon_slave_readdata;
  internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write)))))));
  --assign a2h_avalon_slave_waitrequest_from_sa = a2h_avalon_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_a2h_avalon_slave_waitrequest_from_sa <= a2h_avalon_slave_waitrequest;
  --a2h_avalon_slave_arb_share_counter set values, which is an e_mux
  a2h_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --a2h_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  a2h_avalon_slave_non_bursting_master_requests <= std_logic'('0');
  --a2h_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  a2h_avalon_slave_any_bursting_master_saved_grant <= pcie_to_hibi_4x_sopc_burst_5_downstream_saved_grant_a2h_avalon_slave;
  --a2h_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  a2h_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(a2h_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000") & (a2h_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(a2h_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000") & (a2h_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 11);
  --a2h_avalon_slave_allgrants all slave grants, which is an e_mux
  a2h_avalon_slave_allgrants <= a2h_avalon_slave_grant_vector;
  --a2h_avalon_slave_end_xfer assignment, which is an e_assign
  a2h_avalon_slave_end_xfer <= NOT ((a2h_avalon_slave_waits_for_read OR a2h_avalon_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_a2h_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_a2h_avalon_slave <= a2h_avalon_slave_end_xfer AND (((NOT a2h_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --a2h_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  a2h_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_a2h_avalon_slave AND a2h_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_a2h_avalon_slave AND NOT a2h_avalon_slave_non_bursting_master_requests));
  --a2h_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      a2h_avalon_slave_arb_share_counter <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(a2h_avalon_slave_arb_counter_enable) = '1' then 
        a2h_avalon_slave_arb_share_counter <= a2h_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --a2h_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      a2h_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((a2h_avalon_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_a2h_avalon_slave)) OR ((end_xfer_arb_share_counter_term_a2h_avalon_slave AND NOT a2h_avalon_slave_non_bursting_master_requests)))) = '1' then 
        a2h_avalon_slave_slavearbiterlockenable <= or_reduce(a2h_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_5/downstream a2h/avalon_slave arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_arbiterlock <= a2h_avalon_slave_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_5_downstream_continuerequest;
  --a2h_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  a2h_avalon_slave_slavearbiterlockenable2 <= or_reduce(a2h_avalon_slave_arb_share_counter_next_value);
  --pcie_to_hibi_4x_sopc_burst_5/downstream a2h/avalon_slave arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_arbiterlock2 <= a2h_avalon_slave_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_5_downstream_continuerequest;
  --a2h_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  a2h_avalon_slave_any_continuerequest <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_5_downstream_continuerequest continued request, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_continuerequest <= std_logic'('1');
  internal_pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave AND NOT ((pcie_to_hibi_4x_sopc_burst_5_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave <= (internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave AND pcie_to_hibi_4x_sopc_burst_5_downstream_read) AND NOT a2h_avalon_slave_waits_for_read;
  --a2h_avalon_slave_writedata mux, which is an e_mux
  a2h_avalon_slave_writedata <= pcie_to_hibi_4x_sopc_burst_5_downstream_writedata;
  --master is always granted when requested
  internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave;
  --pcie_to_hibi_4x_sopc_burst_5/downstream saved-grant a2h/avalon_slave, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_saved_grant_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave;
  --allow new arb cycle for a2h/avalon_slave, which is an e_assign
  a2h_avalon_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  a2h_avalon_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  a2h_avalon_slave_master_qreq_vector <= std_logic'('1');
  --a2h_avalon_slave_reset_n assignment, which is an e_assign
  a2h_avalon_slave_reset_n <= reset_n;
  --a2h_avalon_slave_firsttransfer first transaction, which is an e_assign
  a2h_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(a2h_avalon_slave_begins_xfer) = '1'), a2h_avalon_slave_unreg_firsttransfer, a2h_avalon_slave_reg_firsttransfer);
  --a2h_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  a2h_avalon_slave_unreg_firsttransfer <= NOT ((a2h_avalon_slave_slavearbiterlockenable AND a2h_avalon_slave_any_continuerequest));
  --a2h_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      a2h_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(a2h_avalon_slave_begins_xfer) = '1' then 
        a2h_avalon_slave_reg_firsttransfer <= a2h_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --a2h_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  a2h_avalon_slave_beginbursttransfer_internal <= a2h_avalon_slave_begins_xfer;
  --a2h_avalon_slave_read assignment, which is an e_mux
  a2h_avalon_slave_read <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave AND pcie_to_hibi_4x_sopc_burst_5_downstream_read;
  --a2h_avalon_slave_write assignment, which is an e_mux
  a2h_avalon_slave_write <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave AND pcie_to_hibi_4x_sopc_burst_5_downstream_write;
  shifted_address_to_a2h_avalon_slave_from_pcie_to_hibi_4x_sopc_burst_5_downstream <= pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave;
  --a2h_avalon_slave_address mux, which is an e_mux
  a2h_avalon_slave_address <= A_EXT (A_SRL(shifted_address_to_a2h_avalon_slave_from_pcie_to_hibi_4x_sopc_burst_5_downstream,std_logic_vector'("00000000000000000000000000000010")), 23);
  --d1_a2h_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_a2h_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_a2h_avalon_slave_end_xfer <= a2h_avalon_slave_end_xfer;
    end if;

  end process;

  --a2h_avalon_slave_waits_for_read in a cycle, which is an e_mux
  a2h_avalon_slave_waits_for_read <= a2h_avalon_slave_in_a_read_cycle AND internal_a2h_avalon_slave_waitrequest_from_sa;
  --a2h_avalon_slave_in_a_read_cycle assignment, which is an e_assign
  a2h_avalon_slave_in_a_read_cycle <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave AND pcie_to_hibi_4x_sopc_burst_5_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= a2h_avalon_slave_in_a_read_cycle;
  --a2h_avalon_slave_waits_for_write in a cycle, which is an e_mux
  a2h_avalon_slave_waits_for_write <= a2h_avalon_slave_in_a_write_cycle AND internal_a2h_avalon_slave_waitrequest_from_sa;
  --a2h_avalon_slave_in_a_write_cycle assignment, which is an e_assign
  a2h_avalon_slave_in_a_write_cycle <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave AND pcie_to_hibi_4x_sopc_burst_5_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= a2h_avalon_slave_in_a_write_cycle;
  wait_for_a2h_avalon_slave_counter <= std_logic'('0');
  --a2h_avalon_slave_byteenable byte enable port mux, which is an e_mux
  a2h_avalon_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  a2h_avalon_slave_waitrequest_from_sa <= internal_a2h_avalon_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave;
--synthesis translate_off
    --a2h/avalon_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave AND to_std_logic((((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("pcie_to_hibi_4x_sopc_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave a2h/avalon_slave"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("pcie_to_hibi_4x_sopc_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave a2h/avalon_slave"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity dma_control_port_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dma_control_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_control_port_slave_readyfordata : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_dma_control_port_slave_end_xfer : OUT STD_LOGIC;
                 signal dma_control_port_slave_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dma_control_port_slave_chipselect : OUT STD_LOGIC;
                 signal dma_control_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_control_port_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal dma_control_port_slave_reset_n : OUT STD_LOGIC;
                 signal dma_control_port_slave_write_n : OUT STD_LOGIC;
                 signal dma_control_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave : OUT STD_LOGIC
              );
end entity dma_control_port_slave_arbitrator;


architecture europa of dma_control_port_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dma_control_port_slave_allgrants :  STD_LOGIC;
                signal dma_control_port_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal dma_control_port_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal dma_control_port_slave_any_continuerequest :  STD_LOGIC;
                signal dma_control_port_slave_arb_counter_enable :  STD_LOGIC;
                signal dma_control_port_slave_arb_share_counter :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_control_port_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_control_port_slave_arb_share_set_values :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_control_port_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal dma_control_port_slave_begins_xfer :  STD_LOGIC;
                signal dma_control_port_slave_end_xfer :  STD_LOGIC;
                signal dma_control_port_slave_firsttransfer :  STD_LOGIC;
                signal dma_control_port_slave_grant_vector :  STD_LOGIC;
                signal dma_control_port_slave_in_a_read_cycle :  STD_LOGIC;
                signal dma_control_port_slave_in_a_write_cycle :  STD_LOGIC;
                signal dma_control_port_slave_master_qreq_vector :  STD_LOGIC;
                signal dma_control_port_slave_non_bursting_master_requests :  STD_LOGIC;
                signal dma_control_port_slave_reg_firsttransfer :  STD_LOGIC;
                signal dma_control_port_slave_slavearbiterlockenable :  STD_LOGIC;
                signal dma_control_port_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal dma_control_port_slave_unreg_firsttransfer :  STD_LOGIC;
                signal dma_control_port_slave_waits_for_read :  STD_LOGIC;
                signal dma_control_port_slave_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_dma_control_port_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_saved_grant_dma_control_port_slave :  STD_LOGIC;
                signal wait_for_dma_control_port_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT dma_control_port_slave_end_xfer;
    end if;

  end process;

  dma_control_port_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave);
  --assign dma_control_port_slave_readdata_from_sa = dma_control_port_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dma_control_port_slave_readdata_from_sa <= dma_control_port_slave_readdata;
  internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write)))))));
  --assign dma_control_port_slave_readyfordata_from_sa = dma_control_port_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dma_control_port_slave_readyfordata_from_sa <= dma_control_port_slave_readyfordata;
  --dma_control_port_slave_arb_share_counter set values, which is an e_mux
  dma_control_port_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --dma_control_port_slave_non_bursting_master_requests mux, which is an e_mux
  dma_control_port_slave_non_bursting_master_requests <= std_logic'('0');
  --dma_control_port_slave_any_bursting_master_saved_grant mux, which is an e_mux
  dma_control_port_slave_any_bursting_master_saved_grant <= pcie_to_hibi_4x_sopc_burst_4_downstream_saved_grant_dma_control_port_slave;
  --dma_control_port_slave_arb_share_counter_next_value assignment, which is an e_assign
  dma_control_port_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(dma_control_port_slave_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000") & (dma_control_port_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(dma_control_port_slave_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000") & (dma_control_port_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 11);
  --dma_control_port_slave_allgrants all slave grants, which is an e_mux
  dma_control_port_slave_allgrants <= dma_control_port_slave_grant_vector;
  --dma_control_port_slave_end_xfer assignment, which is an e_assign
  dma_control_port_slave_end_xfer <= NOT ((dma_control_port_slave_waits_for_read OR dma_control_port_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_dma_control_port_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_dma_control_port_slave <= dma_control_port_slave_end_xfer AND (((NOT dma_control_port_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --dma_control_port_slave_arb_share_counter arbitration counter enable, which is an e_assign
  dma_control_port_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_dma_control_port_slave AND dma_control_port_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_dma_control_port_slave AND NOT dma_control_port_slave_non_bursting_master_requests));
  --dma_control_port_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_control_port_slave_arb_share_counter <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(dma_control_port_slave_arb_counter_enable) = '1' then 
        dma_control_port_slave_arb_share_counter <= dma_control_port_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --dma_control_port_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_control_port_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((dma_control_port_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_dma_control_port_slave)) OR ((end_xfer_arb_share_counter_term_dma_control_port_slave AND NOT dma_control_port_slave_non_bursting_master_requests)))) = '1' then 
        dma_control_port_slave_slavearbiterlockenable <= or_reduce(dma_control_port_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_4/downstream dma/control_port_slave arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_arbiterlock <= dma_control_port_slave_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_4_downstream_continuerequest;
  --dma_control_port_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  dma_control_port_slave_slavearbiterlockenable2 <= or_reduce(dma_control_port_slave_arb_share_counter_next_value);
  --pcie_to_hibi_4x_sopc_burst_4/downstream dma/control_port_slave arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_arbiterlock2 <= dma_control_port_slave_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_4_downstream_continuerequest;
  --dma_control_port_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  dma_control_port_slave_any_continuerequest <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_4_downstream_continuerequest continued request, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_continuerequest <= std_logic'('1');
  internal_pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave AND NOT ((pcie_to_hibi_4x_sopc_burst_4_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave <= (internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave AND pcie_to_hibi_4x_sopc_burst_4_downstream_read) AND NOT dma_control_port_slave_waits_for_read;
  --dma_control_port_slave_writedata mux, which is an e_mux
  dma_control_port_slave_writedata <= pcie_to_hibi_4x_sopc_burst_4_downstream_writedata;
  --master is always granted when requested
  internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave;
  --pcie_to_hibi_4x_sopc_burst_4/downstream saved-grant dma/control_port_slave, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_saved_grant_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave;
  --allow new arb cycle for dma/control_port_slave, which is an e_assign
  dma_control_port_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  dma_control_port_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  dma_control_port_slave_master_qreq_vector <= std_logic'('1');
  --dma_control_port_slave_reset_n assignment, which is an e_assign
  dma_control_port_slave_reset_n <= reset_n;
  dma_control_port_slave_chipselect <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave;
  --dma_control_port_slave_firsttransfer first transaction, which is an e_assign
  dma_control_port_slave_firsttransfer <= A_WE_StdLogic((std_logic'(dma_control_port_slave_begins_xfer) = '1'), dma_control_port_slave_unreg_firsttransfer, dma_control_port_slave_reg_firsttransfer);
  --dma_control_port_slave_unreg_firsttransfer first transaction, which is an e_assign
  dma_control_port_slave_unreg_firsttransfer <= NOT ((dma_control_port_slave_slavearbiterlockenable AND dma_control_port_slave_any_continuerequest));
  --dma_control_port_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_control_port_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(dma_control_port_slave_begins_xfer) = '1' then 
        dma_control_port_slave_reg_firsttransfer <= dma_control_port_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --dma_control_port_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  dma_control_port_slave_beginbursttransfer_internal <= dma_control_port_slave_begins_xfer;
  --~dma_control_port_slave_write_n assignment, which is an e_mux
  dma_control_port_slave_write_n <= NOT ((internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave AND pcie_to_hibi_4x_sopc_burst_4_downstream_write));
  --dma_control_port_slave_address mux, which is an e_mux
  dma_control_port_slave_address <= pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress (2 DOWNTO 0);
  --d1_dma_control_port_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_dma_control_port_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_dma_control_port_slave_end_xfer <= dma_control_port_slave_end_xfer;
    end if;

  end process;

  --dma_control_port_slave_waits_for_read in a cycle, which is an e_mux
  dma_control_port_slave_waits_for_read <= dma_control_port_slave_in_a_read_cycle AND dma_control_port_slave_begins_xfer;
  --dma_control_port_slave_in_a_read_cycle assignment, which is an e_assign
  dma_control_port_slave_in_a_read_cycle <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave AND pcie_to_hibi_4x_sopc_burst_4_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= dma_control_port_slave_in_a_read_cycle;
  --dma_control_port_slave_waits_for_write in a cycle, which is an e_mux
  dma_control_port_slave_waits_for_write <= dma_control_port_slave_in_a_write_cycle AND dma_control_port_slave_begins_xfer;
  --dma_control_port_slave_in_a_write_cycle assignment, which is an e_assign
  dma_control_port_slave_in_a_write_cycle <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave AND pcie_to_hibi_4x_sopc_burst_4_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= dma_control_port_slave_in_a_write_cycle;
  wait_for_dma_control_port_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave;
--synthesis translate_off
    --dma/control_port_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave AND to_std_logic((((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("pcie_to_hibi_4x_sopc_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave dma/control_port_slave"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("pcie_to_hibi_4x_sopc_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave dma/control_port_slave"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity dma_read_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer : IN STD_LOGIC;
                 signal dma_read_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_read_master_chipselect : IN STD_LOGIC;
                 signal dma_read_master_flush : IN STD_LOGIC;
                 signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                 signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                 signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                 signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal dma_read_master_read_n : IN STD_LOGIC;
                 signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                 signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal dma_read_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_read_master_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dma_read_master_flush_qualified_exported : OUT STD_LOGIC;
                 signal dma_read_master_latency_counter : OUT STD_LOGIC;
                 signal dma_read_master_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal dma_read_master_readdatavalid : OUT STD_LOGIC;
                 signal dma_read_master_waitrequest : OUT STD_LOGIC
              );
end entity dma_read_master_arbitrator;


architecture europa of dma_read_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal dma_read_master_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_read_master_burstcount_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_read_master_chipselect_last_time :  STD_LOGIC;
                signal dma_read_master_dbs_increment :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_read_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_read_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_read_master_flush_qualified :  STD_LOGIC;
                signal dma_read_master_is_granted_some_slave :  STD_LOGIC;
                signal dma_read_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_read_master_read_but_no_slave_selected :  STD_LOGIC;
                signal dma_read_master_read_n_last_time :  STD_LOGIC;
                signal dma_read_master_run :  STD_LOGIC;
                signal dma_read_master_run_delayed :  STD_LOGIC;
                signal internal_dma_read_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_dma_read_master_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_dma_read_master_latency_counter :  STD_LOGIC;
                signal internal_dma_read_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dma_read_master_latency_counter :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_dma_read_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream OR NOT dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream OR NOT dma_read_master_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_read_master_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream OR NOT dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream OR NOT ((NOT dma_read_master_read_n AND dma_read_master_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((NOT dma_read_master_read_n AND dma_read_master_chipselect)))))))))));
  --cascaded wait assignment, which is an e_assign
  dma_read_master_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_dma_read_master_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(dma_read_master_address(31)) & std_logic_vector'("0000000000") & dma_read_master_address(20 DOWNTO 0));
  --dma_read_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_read_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      dma_read_master_read_but_no_slave_selected <= (((NOT dma_read_master_read_n AND dma_read_master_chipselect)) AND dma_read_master_run) AND NOT dma_read_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  dma_read_master_is_granted_some_slave <= dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream OR dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_dma_read_master_readdatavalid <= dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream OR ((dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream AND dbs_rdv_counter_overflow));
  --run delay, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_read_master_run_delayed <= std_logic'('0');
    elsif clk'event and clk = '1' then
      dma_read_master_run_delayed <= dma_read_master_run;
    end if;

  end process;

  --The Flushificator, which is an e_assign
  dma_read_master_flush_qualified <= dma_read_master_flush AND dma_read_master_run_delayed;
  --latent slave read data valid which is not flushed, which is an e_mux
  dma_read_master_readdatavalid <= ((dma_read_master_read_but_no_slave_selected OR ((pre_flush_dma_read_master_readdatavalid AND NOT dma_read_master_flush_qualified))) OR dma_read_master_read_but_no_slave_selected) OR ((pre_flush_dma_read_master_readdatavalid AND NOT dma_read_master_flush_qualified));
  --The Exported Flushificator, which is an e_assign
  dma_read_master_flush_qualified_exported <= dma_read_master_flush_qualified;
  --dma/read_master readdata mux, which is an e_mux
  dma_read_master_readdata <= ((A_REP(NOT dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream, 64) OR pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa)) AND ((A_REP(NOT dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream, 64) OR Std_Logic_Vector'(pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa(31 DOWNTO 0) & dbs_latent_32_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_dma_read_master_waitrequest <= NOT dma_read_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_dma_read_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_dma_read_master_latency_counter <= p1_dma_read_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_dma_read_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((dma_read_master_run AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect))))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_dma_read_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_dma_read_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to latent dbs-32 stored 0, which is an e_mux
  p1_dbs_latent_32_reg_segment_0 <= pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa;
  --dbs register for latent dbs-32 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_0 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((dma_read_master_dbs_rdv_counter(2))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_32_reg_segment_0 <= p1_dbs_latent_32_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  dma_read_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000000")), 3);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_dma_read_master_dbs_address(2) AND NOT((next_dbs_address(2)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_dma_read_master_dbs_address)) + (std_logic_vector'("0") & (dma_read_master_dbs_increment))), 3);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_dma_read_master_dbs_address <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_dma_read_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  dma_read_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (dma_read_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (dma_read_master_dbs_rdv_counter_inc))), 3);
  --dma_read_master_rdv_inc_mux, which is an e_mux
  dma_read_master_dbs_rdv_counter_inc <= std_logic_vector'("100");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dma_read_master_dbs_rdv_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable OR dma_read_master_flush_qualified)) = '1' then 
        if std_logic'(dma_read_master_flush_qualified) = '1' then 
          dma_read_master_dbs_rdv_counter <= std_logic_vector'("000");
        else
          dma_read_master_dbs_rdv_counter <= dma_read_master_next_dbs_rdv_counter;
        end if;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= dma_read_master_dbs_rdv_counter(2) AND NOT dma_read_master_next_dbs_rdv_counter(2);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  dma_read_master_address_to_slave <= internal_dma_read_master_address_to_slave;
  --vhdl renameroo for output signals
  dma_read_master_dbs_address <= internal_dma_read_master_dbs_address;
  --vhdl renameroo for output signals
  dma_read_master_latency_counter <= internal_dma_read_master_latency_counter;
  --vhdl renameroo for output signals
  dma_read_master_waitrequest <= internal_dma_read_master_waitrequest;
--synthesis translate_off
    --dma_read_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_read_master_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        dma_read_master_address_last_time <= dma_read_master_address;
      end if;

    end process;

    --dma/read_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_dma_read_master_waitrequest AND dma_read_master_chipselect;
      end if;

    end process;

    --dma_read_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((dma_read_master_address /= dma_read_master_address_last_time))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("dma_read_master_address did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_read_master_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_read_master_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        dma_read_master_chipselect_last_time <= dma_read_master_chipselect;
      end if;

    end process;

    --dma_read_master_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(dma_read_master_chipselect) /= std_logic'(dma_read_master_chipselect_last_time)))))) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("dma_read_master_chipselect did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_read_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_read_master_burstcount_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        dma_read_master_burstcount_last_time <= dma_read_master_burstcount;
      end if;

    end process;

    --dma_read_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((dma_read_master_burstcount /= dma_read_master_burstcount_last_time))))) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("dma_read_master_burstcount did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --~dma_read_master_read_n check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_read_master_read_n_last_time <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
      elsif clk'event and clk = '1' then
        dma_read_master_read_n_last_time <= dma_read_master_read_n;
      end if;

    end process;

    --~dma_read_master_read_n matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NOT dma_read_master_read_n) /= std_logic'(NOT dma_read_master_read_n_last_time)))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("~dma_read_master_read_n did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity dma_write_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer : IN STD_LOGIC;
                 signal dma_write_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal dma_write_master_chipselect : IN STD_LOGIC;
                 signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                 signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                 signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                 signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                 signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                 signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                 signal dma_write_master_write_n : IN STD_LOGIC;
                 signal dma_write_master_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal dma_write_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dma_write_master_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_waitrequest : OUT STD_LOGIC
              );
end entity dma_write_master_arbitrator;


architecture europa of dma_write_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dma_write_master_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_write_master_burstcount_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_write_master_byteenable_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dma_write_master_chipselect_last_time :  STD_LOGIC;
                signal dma_write_master_dbs_increment :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_write_master_run :  STD_LOGIC;
                signal dma_write_master_write_n_last_time :  STD_LOGIC;
                signal dma_write_master_writedata_last_time :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal internal_dma_write_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_dma_write_master_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_dma_write_master_waitrequest :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream OR NOT dma_write_master_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_write_master_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream OR NOT ((NOT dma_write_master_write_n AND dma_write_master_chipselect)))))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_dma_write_master_dbs_address(2)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((NOT dma_write_master_write_n AND dma_write_master_chipselect)))))))))));
  --cascaded wait assignment, which is an e_assign
  dma_write_master_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_dma_write_master_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(dma_write_master_address(31)) & std_logic_vector'("0000000000") & dma_write_master_address(20 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_dma_write_master_waitrequest <= NOT dma_write_master_run;
  --mux write dbs 1, which is an e_mux
  dma_write_master_dbs_write_32 <= A_WE_StdLogicVector((std_logic'((internal_dma_write_master_dbs_address(2))) = '1'), dma_write_master_writedata(63 DOWNTO 32), dma_write_master_writedata(31 DOWNTO 0));
  --dbs count increment, which is an e_mux
  dma_write_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000000")), 3);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_dma_write_master_dbs_address(2) AND NOT((next_dbs_address(2)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_dma_write_master_dbs_address)) + (std_logic_vector'("0") & (dma_write_master_dbs_increment))), 3);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_dma_write_master_dbs_address <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_dma_write_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  dma_write_master_address_to_slave <= internal_dma_write_master_address_to_slave;
  --vhdl renameroo for output signals
  dma_write_master_dbs_address <= internal_dma_write_master_dbs_address;
  --vhdl renameroo for output signals
  dma_write_master_waitrequest <= internal_dma_write_master_waitrequest;
--synthesis translate_off
    --dma_write_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        dma_write_master_address_last_time <= dma_write_master_address;
      end if;

    end process;

    --dma/write_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_dma_write_master_waitrequest AND dma_write_master_chipselect;
      end if;

    end process;

    --dma_write_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((dma_write_master_address /= dma_write_master_address_last_time))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("dma_write_master_address did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_write_master_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        dma_write_master_chipselect_last_time <= dma_write_master_chipselect;
      end if;

    end process;

    --dma_write_master_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(dma_write_master_chipselect) /= std_logic'(dma_write_master_chipselect_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("dma_write_master_chipselect did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_write_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_burstcount_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        dma_write_master_burstcount_last_time <= dma_write_master_burstcount;
      end if;

    end process;

    --dma_write_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((dma_write_master_burstcount /= dma_write_master_burstcount_last_time))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("dma_write_master_burstcount did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_write_master_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_byteenable_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        dma_write_master_byteenable_last_time <= dma_write_master_byteenable;
      end if;

    end process;

    --dma_write_master_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((dma_write_master_byteenable /= dma_write_master_byteenable_last_time))))) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("dma_write_master_byteenable did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --~dma_write_master_write_n check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_write_n_last_time <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
      elsif clk'event and clk = '1' then
        dma_write_master_write_n_last_time <= dma_write_master_write_n;
      end if;

    end process;

    --~dma_write_master_write_n matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NOT dma_write_master_write_n) /= std_logic'(NOT dma_write_master_write_n_last_time)))))) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("~dma_write_master_write_n did not heed wait!!!"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --dma_write_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        dma_write_master_writedata_last_time <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        dma_write_master_writedata_last_time <= dma_write_master_writedata;
      end if;

    end process;

    --dma_write_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((dma_write_master_writedata /= dma_write_master_writedata_last_time)))) AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect)))) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("dma_write_master_writedata did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_Control_Register_Access_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcie_Control_Register_Access_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Control_Register_Access_waitrequest : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_Control_Register_Access_end_xfer : OUT STD_LOGIC;
                 signal pcie_Control_Register_Access_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal pcie_Control_Register_Access_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_Control_Register_Access_chipselect : OUT STD_LOGIC;
                 signal pcie_Control_Register_Access_read : OUT STD_LOGIC;
                 signal pcie_Control_Register_Access_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Control_Register_Access_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_Control_Register_Access_write : OUT STD_LOGIC;
                 signal pcie_Control_Register_Access_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access : OUT STD_LOGIC
              );
end entity pcie_Control_Register_Access_arbitrator;


architecture europa of pcie_Control_Register_Access_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_Control_Register_Access :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcie_Control_Register_Access_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access :  STD_LOGIC;
                signal last_cycle_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_slave_pcie_Control_Register_Access :  STD_LOGIC;
                signal last_cycle_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_slave_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_Control_Register_Access_allgrants :  STD_LOGIC;
                signal pcie_Control_Register_Access_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_Control_Register_Access_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_Control_Register_Access_any_continuerequest :  STD_LOGIC;
                signal pcie_Control_Register_Access_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_arb_counter_enable :  STD_LOGIC;
                signal pcie_Control_Register_Access_arb_share_counter :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_Control_Register_Access_arb_share_counter_next_value :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_Control_Register_Access_arb_share_set_values :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_Control_Register_Access_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_arbitration_holdoff_internal :  STD_LOGIC;
                signal pcie_Control_Register_Access_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_Control_Register_Access_begins_xfer :  STD_LOGIC;
                signal pcie_Control_Register_Access_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Control_Register_Access_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_end_xfer :  STD_LOGIC;
                signal pcie_Control_Register_Access_firsttransfer :  STD_LOGIC;
                signal pcie_Control_Register_Access_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_in_a_read_cycle :  STD_LOGIC;
                signal pcie_Control_Register_Access_in_a_write_cycle :  STD_LOGIC;
                signal pcie_Control_Register_Access_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_Control_Register_Access_reg_firsttransfer :  STD_LOGIC;
                signal pcie_Control_Register_Access_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Control_Register_Access_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_Control_Register_Access_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_Control_Register_Access_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_Control_Register_Access_waits_for_read :  STD_LOGIC;
                signal pcie_Control_Register_Access_waits_for_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access :  STD_LOGIC;
                signal shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_2_downstream :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_3_downstream :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal wait_for_pcie_Control_Register_Access_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_Control_Register_Access_end_xfer;
    end if;

  end process;

  pcie_Control_Register_Access_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access OR internal_pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access));
  --assign pcie_Control_Register_Access_readdata_from_sa = pcie_Control_Register_Access_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_Control_Register_Access_readdata_from_sa <= pcie_Control_Register_Access_readdata;
  internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write)))))));
  --assign pcie_Control_Register_Access_waitrequest_from_sa = pcie_Control_Register_Access_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_Control_Register_Access_waitrequest_from_sa <= pcie_Control_Register_Access_waitrequest;
  --pcie_Control_Register_Access_arb_share_counter set values, which is an e_mux
  pcie_Control_Register_Access_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 12);
  --pcie_Control_Register_Access_non_bursting_master_requests mux, which is an e_mux
  pcie_Control_Register_Access_non_bursting_master_requests <= std_logic'('0');
  --pcie_Control_Register_Access_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_Control_Register_Access_any_bursting_master_saved_grant <= ((pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access OR pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access) OR pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access) OR pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access;
  --pcie_Control_Register_Access_arb_share_counter_next_value assignment, which is an e_assign
  pcie_Control_Register_Access_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_Control_Register_Access_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_Control_Register_Access_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_Control_Register_Access_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_Control_Register_Access_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 12);
  --pcie_Control_Register_Access_allgrants all slave grants, which is an e_mux
  pcie_Control_Register_Access_allgrants <= (((or_reduce(pcie_Control_Register_Access_grant_vector)) OR (or_reduce(pcie_Control_Register_Access_grant_vector))) OR (or_reduce(pcie_Control_Register_Access_grant_vector))) OR (or_reduce(pcie_Control_Register_Access_grant_vector));
  --pcie_Control_Register_Access_end_xfer assignment, which is an e_assign
  pcie_Control_Register_Access_end_xfer <= NOT ((pcie_Control_Register_Access_waits_for_read OR pcie_Control_Register_Access_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_Control_Register_Access arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_Control_Register_Access <= pcie_Control_Register_Access_end_xfer AND (((NOT pcie_Control_Register_Access_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_Control_Register_Access_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_Control_Register_Access_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_Control_Register_Access AND pcie_Control_Register_Access_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_Control_Register_Access AND NOT pcie_Control_Register_Access_non_bursting_master_requests));
  --pcie_Control_Register_Access_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Control_Register_Access_arb_share_counter <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Control_Register_Access_arb_counter_enable) = '1' then 
        pcie_Control_Register_Access_arb_share_counter <= pcie_Control_Register_Access_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_Control_Register_Access_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Control_Register_Access_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(pcie_Control_Register_Access_master_qreq_vector) AND end_xfer_arb_share_counter_term_pcie_Control_Register_Access)) OR ((end_xfer_arb_share_counter_term_pcie_Control_Register_Access AND NOT pcie_Control_Register_Access_non_bursting_master_requests)))) = '1' then 
        pcie_Control_Register_Access_slavearbiterlockenable <= or_reduce(pcie_Control_Register_Access_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2/downstream pcie/Control_Register_Access arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock <= pcie_Control_Register_Access_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest;
  --pcie_Control_Register_Access_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_Control_Register_Access_slavearbiterlockenable2 <= or_reduce(pcie_Control_Register_Access_arb_share_counter_next_value);
  --pcie_to_hibi_4x_sopc_burst_2/downstream pcie/Control_Register_Access arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock2 <= pcie_Control_Register_Access_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_3/downstream pcie/Control_Register_Access arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock <= pcie_Control_Register_Access_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_3/downstream pcie/Control_Register_Access arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock2 <= pcie_Control_Register_Access_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_3/downstream granted pcie/Control_Register_Access last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_slave_pcie_Control_Register_Access <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_slave_pcie_Control_Register_Access <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Control_Register_Access_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_slave_pcie_Control_Register_Access))))));
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest continued request, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_slave_pcie_Control_Register_Access))) AND std_logic_vector'("00000000000000000000000000000001")));
  --pcie_Control_Register_Access_any_continuerequest at least one master continues requesting, which is an e_mux
  pcie_Control_Register_Access_any_continuerequest <= pcie_to_hibi_4x_sopc_burst_3_downstream_continuerequest OR pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest;
  internal_pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access AND NOT ((((pcie_to_hibi_4x_sopc_burst_2_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock));
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access <= (internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_2_downstream_read) AND NOT pcie_Control_Register_Access_waits_for_read;
  --pcie_Control_Register_Access_writedata mux, which is an e_mux
  pcie_Control_Register_Access_writedata <= A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access)) = '1'), pcie_to_hibi_4x_sopc_burst_2_downstream_writedata, pcie_to_hibi_4x_sopc_burst_3_downstream_writedata);
  internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write)))))));
  --pcie_to_hibi_4x_sopc_burst_2/downstream granted pcie/Control_Register_Access last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_slave_pcie_Control_Register_Access <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_slave_pcie_Control_Register_Access <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Control_Register_Access_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_slave_pcie_Control_Register_Access))))));
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest continued request, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_slave_pcie_Control_Register_Access))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access AND NOT ((((pcie_to_hibi_4x_sopc_burst_3_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock));
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access <= (internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_3_downstream_read) AND NOT pcie_Control_Register_Access_waits_for_read;
  --allow new arb cycle for pcie/Control_Register_Access, which is an e_assign
  pcie_Control_Register_Access_allow_new_arb_cycle <= NOT pcie_to_hibi_4x_sopc_burst_2_downstream_arbiterlock AND NOT pcie_to_hibi_4x_sopc_burst_3_downstream_arbiterlock;
  --pcie_to_hibi_4x_sopc_burst_3/downstream assignment into master qualified-requests vector for pcie/Control_Register_Access, which is an e_assign
  pcie_Control_Register_Access_master_qreq_vector(0) <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access;
  --pcie_to_hibi_4x_sopc_burst_3/downstream grant pcie/Control_Register_Access, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access <= pcie_Control_Register_Access_grant_vector(0);
  --pcie_to_hibi_4x_sopc_burst_3/downstream saved-grant pcie/Control_Register_Access, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access <= pcie_Control_Register_Access_arb_winner(0);
  --pcie_to_hibi_4x_sopc_burst_2/downstream assignment into master qualified-requests vector for pcie/Control_Register_Access, which is an e_assign
  pcie_Control_Register_Access_master_qreq_vector(1) <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access;
  --pcie_to_hibi_4x_sopc_burst_2/downstream grant pcie/Control_Register_Access, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access <= pcie_Control_Register_Access_grant_vector(1);
  --pcie_to_hibi_4x_sopc_burst_2/downstream saved-grant pcie/Control_Register_Access, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access <= pcie_Control_Register_Access_arb_winner(1);
  --pcie/Control_Register_Access chosen-master double-vector, which is an e_assign
  pcie_Control_Register_Access_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((pcie_Control_Register_Access_master_qreq_vector & pcie_Control_Register_Access_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT pcie_Control_Register_Access_master_qreq_vector & NOT pcie_Control_Register_Access_master_qreq_vector))) + (std_logic_vector'("000") & (pcie_Control_Register_Access_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  pcie_Control_Register_Access_arb_winner <= A_WE_StdLogicVector((std_logic'(((pcie_Control_Register_Access_allow_new_arb_cycle AND or_reduce(pcie_Control_Register_Access_grant_vector)))) = '1'), pcie_Control_Register_Access_grant_vector, pcie_Control_Register_Access_saved_chosen_master_vector);
  --saved pcie_Control_Register_Access_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Control_Register_Access_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Control_Register_Access_allow_new_arb_cycle) = '1' then 
        pcie_Control_Register_Access_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(pcie_Control_Register_Access_grant_vector)) = '1'), pcie_Control_Register_Access_grant_vector, pcie_Control_Register_Access_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  pcie_Control_Register_Access_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((pcie_Control_Register_Access_chosen_master_double_vector(1) OR pcie_Control_Register_Access_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((pcie_Control_Register_Access_chosen_master_double_vector(0) OR pcie_Control_Register_Access_chosen_master_double_vector(2)))));
  --pcie/Control_Register_Access chosen master rotated left, which is an e_assign
  pcie_Control_Register_Access_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(pcie_Control_Register_Access_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(pcie_Control_Register_Access_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --pcie/Control_Register_Access's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Control_Register_Access_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(pcie_Control_Register_Access_grant_vector)) = '1' then 
        pcie_Control_Register_Access_arb_addend <= A_WE_StdLogicVector((std_logic'(pcie_Control_Register_Access_end_xfer) = '1'), pcie_Control_Register_Access_chosen_master_rot_left, pcie_Control_Register_Access_grant_vector);
      end if;
    end if;

  end process;

  pcie_Control_Register_Access_chipselect <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access OR internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access;
  --pcie_Control_Register_Access_firsttransfer first transaction, which is an e_assign
  pcie_Control_Register_Access_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_Control_Register_Access_begins_xfer) = '1'), pcie_Control_Register_Access_unreg_firsttransfer, pcie_Control_Register_Access_reg_firsttransfer);
  --pcie_Control_Register_Access_unreg_firsttransfer first transaction, which is an e_assign
  pcie_Control_Register_Access_unreg_firsttransfer <= NOT ((pcie_Control_Register_Access_slavearbiterlockenable AND pcie_Control_Register_Access_any_continuerequest));
  --pcie_Control_Register_Access_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Control_Register_Access_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Control_Register_Access_begins_xfer) = '1' then 
        pcie_Control_Register_Access_reg_firsttransfer <= pcie_Control_Register_Access_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_Control_Register_Access_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_Control_Register_Access_beginbursttransfer_internal <= pcie_Control_Register_Access_begins_xfer;
  --pcie_Control_Register_Access_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  pcie_Control_Register_Access_arbitration_holdoff_internal <= pcie_Control_Register_Access_begins_xfer AND pcie_Control_Register_Access_firsttransfer;
  --pcie_Control_Register_Access_read assignment, which is an e_mux
  pcie_Control_Register_Access_read <= ((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_2_downstream_read)) OR ((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_3_downstream_read));
  --pcie_Control_Register_Access_write assignment, which is an e_mux
  pcie_Control_Register_Access_write <= ((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_2_downstream_write)) OR ((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_3_downstream_write));
  shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_2_downstream <= pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave;
  --pcie_Control_Register_Access_address mux, which is an e_mux
  pcie_Control_Register_Access_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access)) = '1'), (A_SRL(shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_2_downstream,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_3_downstream,std_logic_vector'("00000000000000000000000000000010")))), 12);
  shifted_address_to_pcie_Control_Register_Access_from_pcie_to_hibi_4x_sopc_burst_3_downstream <= pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave;
  --d1_pcie_Control_Register_Access_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_Control_Register_Access_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_Control_Register_Access_end_xfer <= pcie_Control_Register_Access_end_xfer;
    end if;

  end process;

  --pcie_Control_Register_Access_waits_for_read in a cycle, which is an e_mux
  pcie_Control_Register_Access_waits_for_read <= pcie_Control_Register_Access_in_a_read_cycle AND internal_pcie_Control_Register_Access_waitrequest_from_sa;
  --pcie_Control_Register_Access_in_a_read_cycle assignment, which is an e_assign
  pcie_Control_Register_Access_in_a_read_cycle <= ((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_2_downstream_read)) OR ((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_3_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_Control_Register_Access_in_a_read_cycle;
  --pcie_Control_Register_Access_waits_for_write in a cycle, which is an e_mux
  pcie_Control_Register_Access_waits_for_write <= pcie_Control_Register_Access_in_a_write_cycle AND internal_pcie_Control_Register_Access_waitrequest_from_sa;
  --pcie_Control_Register_Access_in_a_write_cycle assignment, which is an e_assign
  pcie_Control_Register_Access_in_a_write_cycle <= ((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_2_downstream_write)) OR ((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access AND pcie_to_hibi_4x_sopc_burst_3_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_Control_Register_Access_in_a_write_cycle;
  wait_for_pcie_Control_Register_Access_counter <= std_logic'('0');
  --pcie_Control_Register_Access_byteenable byte enable port mux, which is an e_mux
  pcie_Control_Register_Access_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  pcie_Control_Register_Access_waitrequest_from_sa <= internal_pcie_Control_Register_Access_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access;
--synthesis translate_off
    --pcie/Control_Register_Access enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access AND to_std_logic((((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("pcie_to_hibi_4x_sopc_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave pcie/Control_Register_Access"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("pcie_to_hibi_4x_sopc_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave pcie/Control_Register_Access"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access AND to_std_logic((((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("pcie_to_hibi_4x_sopc_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave pcie/Control_Register_Access"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("pcie_to_hibi_4x_sopc_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave pcie/Control_Register_Access"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_2_downstream_saved_grant_pcie_Control_Register_Access))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_3_downstream_saved_grant_pcie_Control_Register_Access))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_pcie_Tx_Interface_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_pcie_Tx_Interface_module;


architecture europa of burstcount_fifo_for_pcie_Tx_Interface_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_10 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_11 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_12 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_13 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_14 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_15 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_16 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_17 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_18 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_19 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_20 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_21 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_22 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_23 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_24 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_25 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_26 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_27 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_28 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_29 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_30 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_31 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_9 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic_vector'("0000000000");
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic_vector'("0000000000");
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic_vector'("0000000000");
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic_vector'("0000000000");
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic_vector'("0000000000");
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic_vector'("0000000000");
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic_vector'("0000000000");
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic_vector'("0000000000");
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic_vector'("0000000000");
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic_vector'("0000000000");
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic_vector'("0000000000");
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic_vector'("0000000000");
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic_vector'("0000000000");
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic_vector'("0000000000");
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic_vector'("0000000000");
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic_vector'("0000000000");
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic_vector'("0000000000");
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic_vector'("0000000000");
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic_vector'("0000000000");
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic_vector'("0000000000");
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic_vector'("0000000000");
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic_vector'("0000000000");
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic_vector'("0000000000");
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("0000000000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("0000000000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("0000000000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("0000000000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("0000000000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("0000000000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000000000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module;


architecture europa of rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module;


architecture europa of rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_Tx_Interface_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcie_Tx_Interface_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_Tx_Interface_readdatavalid : IN STD_LOGIC;
                 signal pcie_Tx_Interface_waitrequest : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_Tx_Interface_end_xfer : OUT STD_LOGIC;
                 signal pcie_Tx_Interface_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal pcie_Tx_Interface_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_Tx_Interface_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_Tx_Interface_chipselect : OUT STD_LOGIC;
                 signal pcie_Tx_Interface_read : OUT STD_LOGIC;
                 signal pcie_Tx_Interface_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_Tx_Interface_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_Tx_Interface_write : OUT STD_LOGIC;
                 signal pcie_Tx_Interface_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface : OUT STD_LOGIC
              );
end entity pcie_Tx_Interface_arbitrator;


architecture europa of pcie_Tx_Interface_arbitrator is
component burstcount_fifo_for_pcie_Tx_Interface_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_pcie_Tx_Interface_module;

component rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module;

component rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_Tx_Interface :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcie_Tx_Interface_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_pcie_Tx_Interface_read :  STD_LOGIC;
                signal internal_pcie_Tx_Interface_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_Tx_Interface_write :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface :  STD_LOGIC;
                signal last_cycle_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_slave_pcie_Tx_Interface :  STD_LOGIC;
                signal last_cycle_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_slave_pcie_Tx_Interface :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal p0_pcie_Tx_Interface_load_fifo :  STD_LOGIC;
                signal pcie_Tx_Interface_allgrants :  STD_LOGIC;
                signal pcie_Tx_Interface_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_Tx_Interface_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_Tx_Interface_any_continuerequest :  STD_LOGIC;
                signal pcie_Tx_Interface_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_arb_counter_enable :  STD_LOGIC;
                signal pcie_Tx_Interface_arb_share_counter :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_Tx_Interface_arb_share_counter_next_value :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_Tx_Interface_arb_share_set_values :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_Tx_Interface_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_arbitration_holdoff_internal :  STD_LOGIC;
                signal pcie_Tx_Interface_bbt_burstcounter :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_Tx_Interface_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_Tx_Interface_begins_xfer :  STD_LOGIC;
                signal pcie_Tx_Interface_burstcount_fifo_empty :  STD_LOGIC;
                signal pcie_Tx_Interface_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Tx_Interface_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_current_burst :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_current_burst_minus_one :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_end_xfer :  STD_LOGIC;
                signal pcie_Tx_Interface_firsttransfer :  STD_LOGIC;
                signal pcie_Tx_Interface_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_in_a_read_cycle :  STD_LOGIC;
                signal pcie_Tx_Interface_in_a_write_cycle :  STD_LOGIC;
                signal pcie_Tx_Interface_load_fifo :  STD_LOGIC;
                signal pcie_Tx_Interface_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_move_on_to_next_transaction :  STD_LOGIC;
                signal pcie_Tx_Interface_next_bbt_burstcount :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_Tx_Interface_next_burst_count :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_Tx_Interface_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_Tx_Interface_reg_firsttransfer :  STD_LOGIC;
                signal pcie_Tx_Interface_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcie_Tx_Interface_selected_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_Tx_Interface_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_Tx_Interface_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal pcie_Tx_Interface_transaction_burst_count :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_Tx_Interface_waits_for_read :  STD_LOGIC;
                signal pcie_Tx_Interface_waits_for_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_empty_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_output_from_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_empty_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_output_from_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface :  STD_LOGIC;
                signal shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_0_downstream :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_1_downstream :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal wait_for_pcie_Tx_Interface_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_Tx_Interface_end_xfer;
    end if;

  end process;

  pcie_Tx_Interface_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface OR internal_pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface));
  --assign pcie_Tx_Interface_readdata_from_sa = pcie_Tx_Interface_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_Tx_Interface_readdata_from_sa <= pcie_Tx_Interface_readdata;
  internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write)))))));
  --assign pcie_Tx_Interface_waitrequest_from_sa = pcie_Tx_Interface_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_Tx_Interface_waitrequest_from_sa <= pcie_Tx_Interface_waitrequest;
  --assign pcie_Tx_Interface_readdatavalid_from_sa = pcie_Tx_Interface_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_Tx_Interface_readdatavalid_from_sa <= pcie_Tx_Interface_readdatavalid;
  --pcie_Tx_Interface_arb_share_counter set values, which is an e_mux
  pcie_Tx_Interface_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 11);
  --pcie_Tx_Interface_non_bursting_master_requests mux, which is an e_mux
  pcie_Tx_Interface_non_bursting_master_requests <= std_logic'('0');
  --pcie_Tx_Interface_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_Tx_Interface_any_bursting_master_saved_grant <= ((pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface OR pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface) OR pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface) OR pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface;
  --pcie_Tx_Interface_arb_share_counter_next_value assignment, which is an e_assign
  pcie_Tx_Interface_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_Tx_Interface_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000") & (pcie_Tx_Interface_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_Tx_Interface_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000") & (pcie_Tx_Interface_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 11);
  --pcie_Tx_Interface_allgrants all slave grants, which is an e_mux
  pcie_Tx_Interface_allgrants <= (((or_reduce(pcie_Tx_Interface_grant_vector)) OR (or_reduce(pcie_Tx_Interface_grant_vector))) OR (or_reduce(pcie_Tx_Interface_grant_vector))) OR (or_reduce(pcie_Tx_Interface_grant_vector));
  --pcie_Tx_Interface_end_xfer assignment, which is an e_assign
  pcie_Tx_Interface_end_xfer <= NOT ((pcie_Tx_Interface_waits_for_read OR pcie_Tx_Interface_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_Tx_Interface arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_Tx_Interface <= pcie_Tx_Interface_end_xfer AND (((NOT pcie_Tx_Interface_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_Tx_Interface_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_Tx_Interface_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_Tx_Interface AND pcie_Tx_Interface_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_Tx_Interface AND NOT pcie_Tx_Interface_non_bursting_master_requests));
  --pcie_Tx_Interface_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_arb_share_counter <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Tx_Interface_arb_counter_enable) = '1' then 
        pcie_Tx_Interface_arb_share_counter <= pcie_Tx_Interface_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_Tx_Interface_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(pcie_Tx_Interface_master_qreq_vector) AND end_xfer_arb_share_counter_term_pcie_Tx_Interface)) OR ((end_xfer_arb_share_counter_term_pcie_Tx_Interface AND NOT pcie_Tx_Interface_non_bursting_master_requests)))) = '1' then 
        pcie_Tx_Interface_slavearbiterlockenable <= or_reduce(pcie_Tx_Interface_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0/downstream pcie/Tx_Interface arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock <= pcie_Tx_Interface_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest;
  --pcie_Tx_Interface_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_Tx_Interface_slavearbiterlockenable2 <= or_reduce(pcie_Tx_Interface_arb_share_counter_next_value);
  --pcie_to_hibi_4x_sopc_burst_0/downstream pcie/Tx_Interface arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock2 <= pcie_Tx_Interface_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_1/downstream pcie/Tx_Interface arbiterlock, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock <= pcie_Tx_Interface_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_1/downstream pcie/Tx_Interface arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock2 <= pcie_Tx_Interface_slavearbiterlockenable2 AND pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_1/downstream granted pcie/Tx_Interface last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_slave_pcie_Tx_Interface <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_slave_pcie_Tx_Interface <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Tx_Interface_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_slave_pcie_Tx_Interface))))));
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest continued request, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_slave_pcie_Tx_Interface))) AND std_logic_vector'("00000000000000000000000000000001")));
  --pcie_Tx_Interface_any_continuerequest at least one master continues requesting, which is an e_mux
  pcie_Tx_Interface_any_continuerequest <= pcie_to_hibi_4x_sopc_burst_1_downstream_continuerequest OR pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest;
  internal_pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface AND NOT ((((pcie_to_hibi_4x_sopc_burst_0_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter)))))))))) OR pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock));
  --unique name for pcie_Tx_Interface_move_on_to_next_transaction, which is an e_assign
  pcie_Tx_Interface_move_on_to_next_transaction <= pcie_Tx_Interface_this_cycle_is_the_last_burst AND pcie_Tx_Interface_load_fifo;
  --the currently selected burstcount for pcie_Tx_Interface, which is an e_mux
  pcie_Tx_Interface_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), 10);
  --burstcount_fifo_for_pcie_Tx_Interface, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_pcie_Tx_Interface : burstcount_fifo_for_pcie_Tx_Interface_module
    port map(
      data_out => pcie_Tx_Interface_transaction_burst_count,
      empty => pcie_Tx_Interface_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => pcie_Tx_Interface_selected_burstcount,
      read => pcie_Tx_Interface_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= ((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read) AND pcie_Tx_Interface_load_fifo) AND NOT ((pcie_Tx_Interface_this_cycle_is_the_last_burst AND pcie_Tx_Interface_burstcount_fifo_empty));

  --pcie_Tx_Interface current burst minus one, which is an e_assign
  pcie_Tx_Interface_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000") & (pcie_Tx_Interface_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 10);
  --what to load in current_burst, for pcie_Tx_Interface, which is an e_mux
  pcie_Tx_Interface_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read)) AND NOT pcie_Tx_Interface_load_fifo))) = '1'), pcie_Tx_Interface_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read) AND pcie_Tx_Interface_this_cycle_is_the_last_burst) AND pcie_Tx_Interface_burstcount_fifo_empty))) = '1'), pcie_Tx_Interface_selected_burstcount, A_WE_StdLogicVector((std_logic'((pcie_Tx_Interface_this_cycle_is_the_last_burst)) = '1'), pcie_Tx_Interface_transaction_burst_count, pcie_Tx_Interface_current_burst_minus_one)));
  --the current burst count for pcie_Tx_Interface, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_current_burst <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((pcie_Tx_Interface_readdatavalid_from_sa OR ((NOT pcie_Tx_Interface_load_fifo AND ((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read)))))) = '1' then 
        pcie_Tx_Interface_current_burst <= pcie_Tx_Interface_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_pcie_Tx_Interface_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT pcie_Tx_Interface_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read)) AND pcie_Tx_Interface_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Tx_Interface_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read)) AND NOT pcie_Tx_Interface_load_fifo) OR pcie_Tx_Interface_this_cycle_is_the_last_burst)) = '1' then 
        pcie_Tx_Interface_load_fifo <= p0_pcie_Tx_Interface_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for pcie_Tx_Interface, which is an e_assign
  pcie_Tx_Interface_this_cycle_is_the_last_burst <= NOT (or_reduce(pcie_Tx_Interface_current_burst_minus_one)) AND pcie_Tx_Interface_readdatavalid_from_sa;
  --rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface : rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_0_downstream_to_pcie_Tx_Interface_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_output_from_pcie_Tx_Interface,
      empty => open,
      fifo_contains_ones_n => pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_empty_pcie_Tx_Interface,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface,
      read => pcie_Tx_Interface_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read;

  pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register <= NOT pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_empty_pcie_Tx_Interface;
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface <= ((pcie_Tx_Interface_readdatavalid_from_sa AND pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_output_from_pcie_Tx_Interface)) AND NOT pcie_to_hibi_4x_sopc_burst_0_downstream_rdv_fifo_empty_pcie_Tx_Interface;
  --pcie_Tx_Interface_writedata mux, which is an e_mux
  pcie_Tx_Interface_writedata <= A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), pcie_to_hibi_4x_sopc_burst_0_downstream_writedata, pcie_to_hibi_4x_sopc_burst_1_downstream_writedata);
  internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write)))))));
  --pcie_to_hibi_4x_sopc_burst_0/downstream granted pcie/Tx_Interface last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_slave_pcie_Tx_Interface <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_slave_pcie_Tx_Interface <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Tx_Interface_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_slave_pcie_Tx_Interface))))));
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest continued request, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_slave_pcie_Tx_Interface))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface AND NOT ((((pcie_to_hibi_4x_sopc_burst_1_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter)))))))))) OR pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock));
  --rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface : rdv_fifo_for_pcie_to_hibi_4x_sopc_burst_1_downstream_to_pcie_Tx_Interface_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_output_from_pcie_Tx_Interface,
      empty => open,
      fifo_contains_ones_n => pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_empty_pcie_Tx_Interface,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface,
      read => pcie_Tx_Interface_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT pcie_Tx_Interface_waits_for_read;

  pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register <= NOT pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_empty_pcie_Tx_Interface;
  --local readdatavalid pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface <= ((pcie_Tx_Interface_readdatavalid_from_sa AND pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_output_from_pcie_Tx_Interface)) AND NOT pcie_to_hibi_4x_sopc_burst_1_downstream_rdv_fifo_empty_pcie_Tx_Interface;
  --allow new arb cycle for pcie/Tx_Interface, which is an e_assign
  pcie_Tx_Interface_allow_new_arb_cycle <= NOT pcie_to_hibi_4x_sopc_burst_0_downstream_arbiterlock AND NOT pcie_to_hibi_4x_sopc_burst_1_downstream_arbiterlock;
  --pcie_to_hibi_4x_sopc_burst_1/downstream assignment into master qualified-requests vector for pcie/Tx_Interface, which is an e_assign
  pcie_Tx_Interface_master_qreq_vector(0) <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface;
  --pcie_to_hibi_4x_sopc_burst_1/downstream grant pcie/Tx_Interface, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface <= pcie_Tx_Interface_grant_vector(0);
  --pcie_to_hibi_4x_sopc_burst_1/downstream saved-grant pcie/Tx_Interface, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface <= pcie_Tx_Interface_arb_winner(0);
  --pcie_to_hibi_4x_sopc_burst_0/downstream assignment into master qualified-requests vector for pcie/Tx_Interface, which is an e_assign
  pcie_Tx_Interface_master_qreq_vector(1) <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface;
  --pcie_to_hibi_4x_sopc_burst_0/downstream grant pcie/Tx_Interface, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface <= pcie_Tx_Interface_grant_vector(1);
  --pcie_to_hibi_4x_sopc_burst_0/downstream saved-grant pcie/Tx_Interface, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface <= pcie_Tx_Interface_arb_winner(1);
  --pcie/Tx_Interface chosen-master double-vector, which is an e_assign
  pcie_Tx_Interface_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((pcie_Tx_Interface_master_qreq_vector & pcie_Tx_Interface_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT pcie_Tx_Interface_master_qreq_vector & NOT pcie_Tx_Interface_master_qreq_vector))) + (std_logic_vector'("000") & (pcie_Tx_Interface_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  pcie_Tx_Interface_arb_winner <= A_WE_StdLogicVector((std_logic'(((pcie_Tx_Interface_allow_new_arb_cycle AND or_reduce(pcie_Tx_Interface_grant_vector)))) = '1'), pcie_Tx_Interface_grant_vector, pcie_Tx_Interface_saved_chosen_master_vector);
  --saved pcie_Tx_Interface_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Tx_Interface_allow_new_arb_cycle) = '1' then 
        pcie_Tx_Interface_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(pcie_Tx_Interface_grant_vector)) = '1'), pcie_Tx_Interface_grant_vector, pcie_Tx_Interface_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  pcie_Tx_Interface_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((pcie_Tx_Interface_chosen_master_double_vector(1) OR pcie_Tx_Interface_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((pcie_Tx_Interface_chosen_master_double_vector(0) OR pcie_Tx_Interface_chosen_master_double_vector(2)))));
  --pcie/Tx_Interface chosen master rotated left, which is an e_assign
  pcie_Tx_Interface_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(pcie_Tx_Interface_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(pcie_Tx_Interface_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --pcie/Tx_Interface's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(pcie_Tx_Interface_grant_vector)) = '1' then 
        pcie_Tx_Interface_arb_addend <= A_WE_StdLogicVector((std_logic'(pcie_Tx_Interface_end_xfer) = '1'), pcie_Tx_Interface_chosen_master_rot_left, pcie_Tx_Interface_grant_vector);
      end if;
    end if;

  end process;

  pcie_Tx_Interface_chipselect <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface OR internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface;
  --pcie_Tx_Interface_firsttransfer first transaction, which is an e_assign
  pcie_Tx_Interface_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_Tx_Interface_begins_xfer) = '1'), pcie_Tx_Interface_unreg_firsttransfer, pcie_Tx_Interface_reg_firsttransfer);
  --pcie_Tx_Interface_unreg_firsttransfer first transaction, which is an e_assign
  pcie_Tx_Interface_unreg_firsttransfer <= NOT ((pcie_Tx_Interface_slavearbiterlockenable AND pcie_Tx_Interface_any_continuerequest));
  --pcie_Tx_Interface_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Tx_Interface_begins_xfer) = '1' then 
        pcie_Tx_Interface_reg_firsttransfer <= pcie_Tx_Interface_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_Tx_Interface_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_Tx_Interface_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_Tx_Interface_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_Tx_Interface_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000") & (internal_pcie_Tx_Interface_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_Tx_Interface_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_Tx_Interface_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000") & (pcie_Tx_Interface_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 9);
  --pcie_Tx_Interface_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Tx_Interface_bbt_burstcounter <= std_logic_vector'("000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_Tx_Interface_begins_xfer) = '1' then 
        pcie_Tx_Interface_bbt_burstcounter <= pcie_Tx_Interface_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_Tx_Interface_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_Tx_Interface_beginbursttransfer_internal <= pcie_Tx_Interface_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_Tx_Interface_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_Tx_Interface_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  pcie_Tx_Interface_arbitration_holdoff_internal <= pcie_Tx_Interface_begins_xfer AND pcie_Tx_Interface_firsttransfer;
  --pcie_Tx_Interface_read assignment, which is an e_mux
  internal_pcie_Tx_Interface_read <= ((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_0_downstream_read)) OR ((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_1_downstream_read));
  --pcie_Tx_Interface_write assignment, which is an e_mux
  internal_pcie_Tx_Interface_write <= ((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_0_downstream_write)) OR ((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_1_downstream_write));
  shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_0_downstream <= pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave;
  --pcie_Tx_Interface_address mux, which is an e_mux
  pcie_Tx_Interface_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (A_SRL(shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_0_downstream,std_logic_vector'("00000000000000000000000000000011"))), (A_SRL(shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_1_downstream,std_logic_vector'("00000000000000000000000000000011")))), 18);
  shifted_address_to_pcie_Tx_Interface_from_pcie_to_hibi_4x_sopc_burst_1_downstream <= pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave;
  --d1_pcie_Tx_Interface_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_Tx_Interface_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_Tx_Interface_end_xfer <= pcie_Tx_Interface_end_xfer;
    end if;

  end process;

  --pcie_Tx_Interface_waits_for_read in a cycle, which is an e_mux
  pcie_Tx_Interface_waits_for_read <= pcie_Tx_Interface_in_a_read_cycle AND internal_pcie_Tx_Interface_waitrequest_from_sa;
  --pcie_Tx_Interface_in_a_read_cycle assignment, which is an e_assign
  pcie_Tx_Interface_in_a_read_cycle <= ((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_0_downstream_read)) OR ((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_1_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_Tx_Interface_in_a_read_cycle;
  --pcie_Tx_Interface_waits_for_write in a cycle, which is an e_mux
  pcie_Tx_Interface_waits_for_write <= pcie_Tx_Interface_in_a_write_cycle AND internal_pcie_Tx_Interface_waitrequest_from_sa;
  --pcie_Tx_Interface_in_a_write_cycle assignment, which is an e_assign
  pcie_Tx_Interface_in_a_write_cycle <= ((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_0_downstream_write)) OR ((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface AND pcie_to_hibi_4x_sopc_burst_1_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_Tx_Interface_in_a_write_cycle;
  wait_for_pcie_Tx_Interface_counter <= std_logic'('0');
  --pcie_Tx_Interface_byteenable byte enable port mux, which is an e_mux
  pcie_Tx_Interface_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 8);
  --burstcount mux, which is an e_mux
  internal_pcie_Tx_Interface_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount)), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), 10);
  --vhdl renameroo for output signals
  pcie_Tx_Interface_burstcount <= internal_pcie_Tx_Interface_burstcount;
  --vhdl renameroo for output signals
  pcie_Tx_Interface_read <= internal_pcie_Tx_Interface_read;
  --vhdl renameroo for output signals
  pcie_Tx_Interface_waitrequest_from_sa <= internal_pcie_Tx_Interface_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_Tx_Interface_write <= internal_pcie_Tx_Interface_write;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface;
--synthesis translate_off
    --pcie/Tx_Interface enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface AND to_std_logic((((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("pcie_to_hibi_4x_sopc_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave pcie/Tx_Interface"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("pcie_to_hibi_4x_sopc_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave pcie/Tx_Interface"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface AND to_std_logic((((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("pcie_to_hibi_4x_sopc_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave pcie/Tx_Interface"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("pcie_to_hibi_4x_sopc_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave pcie/Tx_Interface"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_0_downstream_saved_grant_pcie_Tx_Interface))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_1_downstream_saved_grant_pcie_Tx_Interface))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_Rx_Interface_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer : IN STD_LOGIC;
                 signal pcie_Rx_Interface_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                 signal pcie_Rx_Interface_write : IN STD_LOGIC;
                 signal pcie_Rx_Interface_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_Rx_Interface_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pcie_Rx_Interface_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_latency_counter : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_Rx_Interface_readdatavalid : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_reset_n : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_waitrequest : OUT STD_LOGIC
              );
end entity pcie_Rx_Interface_arbitrator;


architecture europa of pcie_Rx_Interface_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_pcie_Rx_Interface_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_pcie_Rx_Interface_latency_counter :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_pcie_Rx_Interface_latency_counter :  STD_LOGIC;
                signal pcie_Rx_Interface_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Rx_Interface_burstcount_last_time :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Rx_Interface_byteenable_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_Rx_Interface_dbs_increment :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pcie_Rx_Interface_dbs_rdv_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pcie_Rx_Interface_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pcie_Rx_Interface_is_granted_some_slave :  STD_LOGIC;
                signal pcie_Rx_Interface_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pcie_Rx_Interface_read_but_no_slave_selected :  STD_LOGIC;
                signal pcie_Rx_Interface_read_last_time :  STD_LOGIC;
                signal pcie_Rx_Interface_run :  STD_LOGIC;
                signal pcie_Rx_Interface_write_last_time :  STD_LOGIC;
                signal pcie_Rx_Interface_writedata_last_time :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_pcie_Rx_Interface_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream OR NOT pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream OR NOT ((pcie_Rx_Interface_read OR pcie_Rx_Interface_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_Rx_Interface_read OR pcie_Rx_Interface_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream OR NOT ((pcie_Rx_Interface_read OR pcie_Rx_Interface_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_Rx_Interface_read OR pcie_Rx_Interface_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream OR NOT pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream OR NOT pcie_Rx_Interface_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream OR NOT pcie_Rx_Interface_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcie_Rx_Interface_dbs_address(2)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_write)))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_Rx_Interface_run <= r_0;
  --pcie_Rx_Interface_reset_n assignment, which is an e_assign
  pcie_Rx_Interface_reset_n <= reset_n;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_Rx_Interface_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(pcie_Rx_Interface_address(31)) & std_logic_vector'("000000") & pcie_Rx_Interface_address(24 DOWNTO 0));
  --pcie_Rx_Interface_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Rx_Interface_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcie_Rx_Interface_read_but_no_slave_selected <= (pcie_Rx_Interface_read AND pcie_Rx_Interface_run) AND NOT pcie_Rx_Interface_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcie_Rx_Interface_is_granted_some_slave <= pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream OR pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_Rx_Interface_readdatavalid <= pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream OR ((pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream AND dbs_rdv_counter_overflow));
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_Rx_Interface_readdatavalid <= ((pcie_Rx_Interface_read_but_no_slave_selected OR pre_flush_pcie_Rx_Interface_readdatavalid) OR pcie_Rx_Interface_read_but_no_slave_selected) OR pre_flush_pcie_Rx_Interface_readdatavalid;
  --pcie/Rx_Interface readdata mux, which is an e_mux
  pcie_Rx_Interface_readdata <= ((A_REP(NOT pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream, 64) OR (std_logic_vector'("00000000000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa)))) AND ((A_REP(NOT pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream, 64) OR Std_Logic_Vector'(pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa(31 DOWNTO 0) & dbs_latent_32_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_pcie_Rx_Interface_waitrequest <= NOT pcie_Rx_Interface_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_Rx_Interface_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcie_Rx_Interface_latency_counter <= p1_pcie_Rx_Interface_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcie_Rx_Interface_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pcie_Rx_Interface_run AND pcie_Rx_Interface_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pcie_Rx_Interface_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to latent dbs-32 stored 0, which is an e_mux
  p1_dbs_latent_32_reg_segment_0 <= pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa;
  --dbs register for latent dbs-32 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_0 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcie_Rx_Interface_dbs_rdv_counter(2))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_32_reg_segment_0 <= p1_dbs_latent_32_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  pcie_Rx_Interface_dbs_write_32 <= A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_dbs_address(2))) = '1'), pcie_Rx_Interface_writedata(63 DOWNTO 32), pcie_Rx_Interface_writedata(31 DOWNTO 0));
  --dbs count increment, which is an e_mux
  pcie_Rx_Interface_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000000")), 3);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_pcie_Rx_Interface_dbs_address(2) AND NOT((next_dbs_address(2)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_pcie_Rx_Interface_dbs_address)) + (std_logic_vector'("0") & (pcie_Rx_Interface_dbs_increment))), 3);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_Rx_Interface_dbs_address <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_pcie_Rx_Interface_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  pcie_Rx_Interface_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (pcie_Rx_Interface_dbs_rdv_counter)) + (std_logic_vector'("0") & (pcie_Rx_Interface_dbs_rdv_counter_inc))), 3);
  --pcie_Rx_Interface_rdv_inc_mux, which is an e_mux
  pcie_Rx_Interface_dbs_rdv_counter_inc <= std_logic_vector'("100");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_Rx_Interface_dbs_rdv_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        pcie_Rx_Interface_dbs_rdv_counter <= pcie_Rx_Interface_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= pcie_Rx_Interface_dbs_rdv_counter(2) AND NOT pcie_Rx_Interface_next_dbs_rdv_counter(2);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa)))))));
  --vhdl renameroo for output signals
  pcie_Rx_Interface_address_to_slave <= internal_pcie_Rx_Interface_address_to_slave;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_dbs_address <= internal_pcie_Rx_Interface_dbs_address;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_latency_counter <= internal_pcie_Rx_Interface_latency_counter;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_waitrequest <= internal_pcie_Rx_Interface_waitrequest;
--synthesis translate_off
    --pcie_Rx_Interface_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_address_last_time <= pcie_Rx_Interface_address;
      end if;

    end process;

    --pcie/Rx_Interface waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_Rx_Interface_waitrequest AND ((pcie_Rx_Interface_read OR pcie_Rx_Interface_write));
      end if;

    end process;

    --pcie_Rx_Interface_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_Rx_Interface_address /= pcie_Rx_Interface_address_last_time))))) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("pcie_Rx_Interface_address did not heed wait!!!"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_Rx_Interface_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_burstcount_last_time <= std_logic_vector'("0000000000");
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_burstcount_last_time <= pcie_Rx_Interface_burstcount;
      end if;

    end process;

    --pcie_Rx_Interface_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_Rx_Interface_burstcount /= pcie_Rx_Interface_burstcount_last_time))))) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("pcie_Rx_Interface_burstcount did not heed wait!!!"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_Rx_Interface_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_byteenable_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_byteenable_last_time <= pcie_Rx_Interface_byteenable;
      end if;

    end process;

    --pcie_Rx_Interface_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_Rx_Interface_byteenable /= pcie_Rx_Interface_byteenable_last_time))))) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("pcie_Rx_Interface_byteenable did not heed wait!!!"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_Rx_Interface_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_read_last_time <= pcie_Rx_Interface_read;
      end if;

    end process;

    --pcie_Rx_Interface_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_Rx_Interface_read) /= std_logic'(pcie_Rx_Interface_read_last_time)))))) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("pcie_Rx_Interface_read did not heed wait!!!"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_Rx_Interface_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_write_last_time <= pcie_Rx_Interface_write;
      end if;

    end process;

    --pcie_Rx_Interface_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_Rx_Interface_write) /= std_logic'(pcie_Rx_Interface_write_last_time)))))) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("pcie_Rx_Interface_write did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_Rx_Interface_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_Rx_Interface_writedata_last_time <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_Rx_Interface_writedata_last_time <= pcie_Rx_Interface_writedata;
      end if;

    end process;

    --pcie_Rx_Interface_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_Rx_Interface_writedata /= pcie_Rx_Interface_writedata_last_time)))) AND pcie_Rx_Interface_write)) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("pcie_Rx_Interface_writedata did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module;


architecture europa of burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_10 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_11 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_12 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_13 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_14 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_15 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_16 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_17 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_18 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_19 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_20 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_21 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_22 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_23 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_24 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_25 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_26 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_27 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_28 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_29 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_30 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_31 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_32 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_33 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_9 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_33;
  empty <= NOT(full_0);
  full_34 <= std_logic'('0');
  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic_vector'("00000000000");
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic_vector'("00000000000");
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic_vector'("00000000000");
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic_vector'("00000000000");
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic_vector'("00000000000");
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic_vector'("00000000000");
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic_vector'("00000000000");
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic_vector'("00000000000");
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic_vector'("00000000000");
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic_vector'("00000000000");
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic_vector'("00000000000");
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic_vector'("00000000000");
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic_vector'("00000000000");
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic_vector'("00000000000");
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic_vector'("00000000000");
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic_vector'("00000000000");
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic_vector'("00000000000");
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic_vector'("00000000000");
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic_vector'("00000000000");
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic_vector'("00000000000");
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic_vector'("00000000000");
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic_vector'("00000000000");
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic_vector'("00000000000");
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic_vector'("00000000000");
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic_vector'("00000000000");
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000000000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000000000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000000000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000000000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000000000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000000000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000000000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module;


architecture europa of rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_33;
  empty <= NOT(full_0);
  full_34 <= std_logic'('0');
  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dma_read_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_read_master_chipselect : IN STD_LOGIC;
                 signal dma_read_master_flush_qualified_exported : IN STD_LOGIC;
                 signal dma_read_master_latency_counter : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal dma_read_master_read_n : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                 signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                 signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : OUT STD_LOGIC;
                 signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_upstream_write : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator is
component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module;

component rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dma_read_master_arbiterlock :  STD_LOGIC;
                signal dma_read_master_arbiterlock2 :  STD_LOGIC;
                signal dma_read_master_continuerequest :  STD_LOGIC;
                signal dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_0_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_upstream_write :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal p0_pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_next_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_selected_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_write :  STD_LOGIC;
                signal wait_for_pcie_to_hibi_4x_sopc_burst_0_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_0_upstream_readdata;
  internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream <= ((to_std_logic(((Std_Logic_Vector'(dma_read_master_address_to_slave(31 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND dma_read_master_chipselect)) AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --assign pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest;
  --assign pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_set_values <= std_logic_vector'("0000000000001");
  --pcie_to_hibi_4x_sopc_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_any_bursting_master_saved_grant <= dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_0_upstream_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 13);
  --pcie_to_hibi_4x_sopc_burst_0_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_0_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream <= pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_0_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream AND pcie_to_hibi_4x_sopc_burst_0_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter <= std_logic_vector'("0000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_0_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_0_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_0_upstream AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --dma/read_master pcie_to_hibi_4x_sopc_burst_0/upstream arbiterlock, which is an e_assign
  dma_read_master_arbiterlock <= pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable AND dma_read_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_0_upstream_arb_share_counter_next_value);
  --dma/read_master pcie_to_hibi_4x_sopc_burst_0/upstream arbiterlock2, which is an e_assign
  dma_read_master_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable2 AND dma_read_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_any_continuerequest <= std_logic'('1');
  --dma_read_master_continuerequest continued request, which is an e_assign
  dma_read_master_continuerequest <= std_logic'('1');
  internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream AND NOT ((((NOT dma_read_master_read_n AND dma_read_master_chipselect)) AND ((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_read_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_read_master_latency_counter))))))) OR (dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register)))));
  --unique name for pcie_to_hibi_4x_sopc_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_move_on_to_next_transaction <= pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo;
  --the currently selected burstcount for pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream : burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_0_upstream_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_0_upstream_transaction_burst_count,
      empty => pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => pcie_to_hibi_4x_sopc_burst_0_upstream_selected_burstcount,
      read => pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo) AND NOT ((pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount_fifo_empty));

  --pcie_to_hibi_4x_sopc_burst_0_upstream current burst minus one, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 11);
  --what to load in current_burst, for pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo))) = '1'), pcie_to_hibi_4x_sopc_burst_0_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst) AND pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount_fifo_empty))) = '1'), pcie_to_hibi_4x_sopc_burst_0_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst)) = '1'), pcie_to_hibi_4x_sopc_burst_0_upstream_transaction_burst_count, pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst_minus_one)));
  --the current burst count for pcie_to_hibi_4x_sopc_burst_0_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa OR ((NOT pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo AND ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read)))))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst <= pcie_to_hibi_4x_sopc_burst_0_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read)) AND pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo) OR pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst)) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo <= p0_pcie_to_hibi_4x_sopc_burst_0_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(pcie_to_hibi_4x_sopc_burst_0_upstream_current_burst_minus_one)) AND pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream : rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_0_upstream_module
    port map(
      data_out => dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_0_upstream,
      empty => open,
      fifo_contains_ones_n => dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_0_upstream,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream,
      read => pcie_to_hibi_4x_sopc_burst_0_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => dma_read_master_flush_qualified_exported,
      write => module_input13
    );

  module_input12 <= std_logic'('0');
  module_input13 <= in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read;

  dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register <= NOT dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --local readdatavalid dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_mux
  dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream <= ((pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid_from_sa AND dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_0_upstream)) AND NOT dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_0/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress <= dma_read_master_address_to_slave (23 DOWNTO 0);
  --master is always granted when requested
  internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --dma/read_master saved-grant pcie_to_hibi_4x_sopc_burst_0/upstream, which is an e_assign
  dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_0/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_0_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_0_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_0_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_0_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_0_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_0_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_0_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_0_upstream_write) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("0000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_0_upstream_read) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 10);
  --pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_0_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_0_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_0_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_0_upstream_read <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --pcie_to_hibi_4x_sopc_burst_0_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_0_upstream_write <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_0_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_address <= dma_read_master_address_to_slave (20 DOWNTO 0);
  --d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_read_cycle <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_0_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_0_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 8);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --vhdl renameroo for output signals
  dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --vhdl renameroo for output signals
  dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_0_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_0_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_0/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --dma/read_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream AND to_std_logic((((std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("dma/read_master drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_0/upstream"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_Tx_Interface_end_xfer : IN STD_LOGIC;
                 signal pcie_Tx_Interface_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_Tx_Interface_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_address : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_last_time :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount_last_time :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_is_granted_some_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata_last_time :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface OR NOT pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface OR NOT pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface OR NOT ((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Tx_Interface_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface OR NOT ((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Tx_Interface_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_0_downstream_address;
  --pcie_to_hibi_4x_sopc_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_but_no_slave_selected <= (pcie_to_hibi_4x_sopc_burst_0_downstream_read AND pcie_to_hibi_4x_sopc_burst_0_downstream_run) AND NOT pcie_to_hibi_4x_sopc_burst_0_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_downstream_is_granted_some_slave <= pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid <= pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface;
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid <= pcie_to_hibi_4x_sopc_burst_0_downstream_read_but_no_slave_selected OR pre_flush_pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_0/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_0_downstream_readdata <= pcie_Tx_Interface_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_0_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter <= p1_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pcie_to_hibi_4x_sopc_burst_0_downstream_run AND pcie_to_hibi_4x_sopc_burst_0_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_0_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_address_last_time <= std_logic_vector'("000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_0_downstream_read OR pcie_to_hibi_4x_sopc_burst_0_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_0_downstream_address /= pcie_to_hibi_4x_sopc_burst_0_downstream_address_last_time))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_address did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount_last_time <= std_logic_vector'("0000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount /= pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount_last_time))))) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable_last_time))))) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_0_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_0_downstream_read_last_time)))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_read did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_0_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_0_downstream_write_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_write did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_writedata_last_time <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_0_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_0_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_0_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_0_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_0_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_0_downstream_write)) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("pcie_to_hibi_4x_sopc_burst_0_downstream_writedata did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dma_write_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal dma_write_master_chipselect : IN STD_LOGIC;
                 signal dma_write_master_write_n : IN STD_LOGIC;
                 signal dma_write_master_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                 signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                 signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                 signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_write : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_upstream_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
              );
end entity pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dma_write_master_arbiterlock :  STD_LOGIC;
                signal dma_write_master_arbiterlock2 :  STD_LOGIC;
                signal dma_write_master_continuerequest :  STD_LOGIC;
                signal dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_1_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_write :  STD_LOGIC;
                signal wait_for_pcie_to_hibi_4x_sopc_burst_1_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_1_upstream_readdata;
  internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream <= ((to_std_logic(((Std_Logic_Vector'(dma_write_master_address_to_slave(31 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND dma_write_master_chipselect)) AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --assign pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_write_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 13);
  --pcie_to_hibi_4x_sopc_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_any_bursting_master_saved_grant <= dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_1_upstream_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 13);
  --pcie_to_hibi_4x_sopc_burst_1_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_1_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream <= pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_1_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream AND pcie_to_hibi_4x_sopc_burst_1_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream AND NOT pcie_to_hibi_4x_sopc_burst_1_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter <= std_logic_vector'("0000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_1_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_1_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_1_upstream AND NOT pcie_to_hibi_4x_sopc_burst_1_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --dma/write_master pcie_to_hibi_4x_sopc_burst_1/upstream arbiterlock, which is an e_assign
  dma_write_master_arbiterlock <= pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable AND dma_write_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_1_upstream_arb_share_counter_next_value);
  --dma/write_master pcie_to_hibi_4x_sopc_burst_1/upstream arbiterlock2, which is an e_assign
  dma_write_master_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable2 AND dma_write_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_any_continuerequest <= std_logic'('1');
  --dma_write_master_continuerequest continued request, which is an e_assign
  dma_write_master_continuerequest <= std_logic'('1');
  internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_writedata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_writedata <= dma_write_master_writedata;
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_1/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress <= dma_write_master_address_to_slave (23 DOWNTO 0);
  --master is always granted when requested
  internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --dma/write_master saved-grant pcie_to_hibi_4x_sopc_burst_1/upstream, which is an e_assign
  dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_1/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_1_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_1_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_1_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_1_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_1_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_1_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_1_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_1_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_1_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_1_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_1_upstream_write) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("0000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_1_upstream_read) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 10);
  --pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_1_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_1_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_1_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_1_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_1_upstream_read <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_1_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_1_upstream_write <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --pcie_to_hibi_4x_sopc_burst_1_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_address <= dma_write_master_address_to_slave (20 DOWNTO 0);
  --d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_read_cycle <= std_logic'('0');
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa;
  --assign pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_write_cycle <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_1_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_1_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream)) = '1'), (std_logic_vector'("000000000000000000000000") & (dma_write_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 8);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_write_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --vhdl renameroo for output signals
  dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --vhdl renameroo for output signals
  dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_1_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_1_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_1/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --dma/write_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream AND to_std_logic((((std_logic_vector'("000000000000000000000") & (dma_write_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("dma/write_master drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_1/upstream"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_Tx_Interface_end_xfer : IN STD_LOGIC;
                 signal pcie_Tx_Interface_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_Tx_Interface_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_address : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_last_time :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount_last_time :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_is_granted_some_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata_last_time :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface OR NOT pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface OR NOT pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface OR NOT ((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Tx_Interface_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface OR NOT ((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Tx_Interface_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_1_downstream_address;
  --pcie_to_hibi_4x_sopc_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_but_no_slave_selected <= (pcie_to_hibi_4x_sopc_burst_1_downstream_read AND pcie_to_hibi_4x_sopc_burst_1_downstream_run) AND NOT pcie_to_hibi_4x_sopc_burst_1_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_downstream_is_granted_some_slave <= pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid <= pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface;
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid <= pcie_to_hibi_4x_sopc_burst_1_downstream_read_but_no_slave_selected OR pre_flush_pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_1/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_1_downstream_readdata <= pcie_Tx_Interface_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_1_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter <= p1_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pcie_to_hibi_4x_sopc_burst_1_downstream_run AND pcie_to_hibi_4x_sopc_burst_1_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_1_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_address_last_time <= std_logic_vector'("000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_1_downstream_read OR pcie_to_hibi_4x_sopc_burst_1_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_1_downstream_address /= pcie_to_hibi_4x_sopc_burst_1_downstream_address_last_time))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_address did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount_last_time <= std_logic_vector'("0000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount /= pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount_last_time))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable_last_time))))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_1_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_1_downstream_read_last_time)))))) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_read did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_1_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_1_downstream_write_last_time)))))) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_write did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_writedata_last_time <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_1_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_1_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_1_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_1_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_1_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_1_downstream_write)) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("pcie_to_hibi_4x_sopc_burst_1_downstream_writedata did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dma_write_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal dma_write_master_chipselect : IN STD_LOGIC;
                 signal dma_write_master_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dma_write_master_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_write_master_write_n : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                 signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                 signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                 signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_write : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dma_write_master_arbiterlock :  STD_LOGIC;
                signal dma_write_master_arbiterlock2 :  STD_LOGIC;
                signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal dma_write_master_continuerequest :  STD_LOGIC;
                signal dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_2_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_write :  STD_LOGIC;
                signal wait_for_pcie_to_hibi_4x_sopc_burst_2_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_2_upstream_readdata;
  internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream <= ((to_std_logic(((Std_Logic_Vector'(dma_write_master_address_to_slave(31 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("10000000000000000100000000000000")))) AND dma_write_master_chipselect)) AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --assign pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & ((A_SLL(dma_write_master_burstcount,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 13);
  --pcie_to_hibi_4x_sopc_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_any_bursting_master_saved_grant <= dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_2_upstream_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 13);
  --pcie_to_hibi_4x_sopc_burst_2_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_2_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream <= pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_2_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream AND pcie_to_hibi_4x_sopc_burst_2_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream AND NOT pcie_to_hibi_4x_sopc_burst_2_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter <= std_logic_vector'("0000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_2_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_2_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_2_upstream AND NOT pcie_to_hibi_4x_sopc_burst_2_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --dma/write_master pcie_to_hibi_4x_sopc_burst_2/upstream arbiterlock, which is an e_assign
  dma_write_master_arbiterlock <= pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable AND dma_write_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_2_upstream_arb_share_counter_next_value);
  --dma/write_master pcie_to_hibi_4x_sopc_burst_2/upstream arbiterlock2, which is an e_assign
  dma_write_master_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable2 AND dma_write_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_any_continuerequest <= std_logic'('1');
  --dma_write_master_continuerequest continued request, which is an e_assign
  dma_write_master_continuerequest <= std_logic'('1');
  internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_writedata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_writedata <= dma_write_master_dbs_write_32;
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_2/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress <= dma_write_master_address_to_slave (15 DOWNTO 0);
  --master is always granted when requested
  internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --dma/write_master saved-grant pcie_to_hibi_4x_sopc_burst_2/upstream, which is an e_assign
  dma_write_master_saved_grant_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_2/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_2_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_2_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_2_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_2_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_2_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_2_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_2_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_2_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_2_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_2_upstream_write) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("0000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_2_upstream_read) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 10);
  --pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_2_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_2_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_2_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_2_upstream_read <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_2_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_2_upstream_write <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --assign pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(dma_write_master_address_to_slave,std_logic_vector'("00000000000000000000000000000011")) & A_ToStdLogicVector(dma_write_master_dbs_address(2)) & A_REP(std_logic'('0'), 2)), 14);
  --d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_read_cycle <= std_logic'('0');
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_write_cycle <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream AND ((NOT dma_write_master_write_n AND dma_write_master_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_2_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_2_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (internal_dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  (dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1(3), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1(2), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1(1), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1(0), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0(3), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0(2), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0(1), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0(0)) <= dma_write_master_byteenable;
  internal_dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_write_master_dbs_address(2)))) = std_logic_vector'("00000000000000000000000000000000"))), dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_0, dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream_segment_1);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_write_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --vhdl renameroo for output signals
  dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --vhdl renameroo for output signals
  dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --vhdl renameroo for output signals
  dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream <= internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_2_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_2_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_2/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --dma/write_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream AND to_std_logic((((std_logic_vector'("000000000000000000000") & (dma_write_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("dma/write_master drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_2/upstream"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_Control_Register_Access_end_xfer : IN STD_LOGIC;
                 signal pcie_Control_Register_Access_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Control_Register_Access_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_last_time :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_is_granted_some_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access OR NOT pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access OR NOT pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access OR NOT ((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Control_Register_Access_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access OR NOT ((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Control_Register_Access_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_2_downstream_address;
  --pcie_to_hibi_4x_sopc_burst_2_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_2_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcie_to_hibi_4x_sopc_burst_2_downstream_read_but_no_slave_selected <= (pcie_to_hibi_4x_sopc_burst_2_downstream_read AND pcie_to_hibi_4x_sopc_burst_2_downstream_run) AND NOT pcie_to_hibi_4x_sopc_burst_2_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_downstream_is_granted_some_slave <= pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid <= (pcie_to_hibi_4x_sopc_burst_2_downstream_read_but_no_slave_selected OR pre_flush_pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid) OR pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access;
  --pcie_to_hibi_4x_sopc_burst_2/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_2_downstream_readdata <= pcie_Control_Register_Access_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_2_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter <= p1_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pcie_to_hibi_4x_sopc_burst_2_downstream_run AND pcie_to_hibi_4x_sopc_burst_2_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_2_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_address_last_time <= std_logic_vector'("00000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_2_downstream_read OR pcie_to_hibi_4x_sopc_burst_2_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_2_downstream_address /= pcie_to_hibi_4x_sopc_burst_2_downstream_address_last_time))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_address did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount) /= std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable_last_time))))) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_read_last_time)))))) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_read did not heed wait!!!"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_2_downstream_write_last_time)))))) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_write did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_2_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_2_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_2_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_2_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_2_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_2_downstream_write)) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("pcie_to_hibi_4x_sopc_burst_2_downstream_writedata did not heed wait!!!"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module;


architecture europa of burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module;


architecture europa of rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dma_read_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal dma_read_master_chipselect : IN STD_LOGIC;
                 signal dma_read_master_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dma_read_master_flush_qualified_exported : IN STD_LOGIC;
                 signal dma_read_master_latency_counter : IN STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal dma_read_master_read_n : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                 signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                 signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                 signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : OUT STD_LOGIC;
                 signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_upstream_write : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator is
component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module;

component rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dma_read_master_arbiterlock :  STD_LOGIC;
                signal dma_read_master_arbiterlock2 :  STD_LOGIC;
                signal dma_read_master_continuerequest :  STD_LOGIC;
                signal dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_3_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_upstream_write :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal p0_pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_next_burst_count :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_selected_burstcount :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_write :  STD_LOGIC;
                signal wait_for_pcie_to_hibi_4x_sopc_burst_3_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid;
  --assign pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_3_upstream_readdata;
  internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream <= ((to_std_logic(((Std_Logic_Vector'(dma_read_master_address_to_slave(31 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("10000000000000000100000000000000")))) AND dma_read_master_chipselect)) AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --assign pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_set_values <= std_logic_vector'("0000000000001");
  --pcie_to_hibi_4x_sopc_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_any_bursting_master_saved_grant <= dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_3_upstream_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 13);
  --pcie_to_hibi_4x_sopc_burst_3_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_3_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream <= pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_3_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream AND pcie_to_hibi_4x_sopc_burst_3_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter <= std_logic_vector'("0000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_3_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_3_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_3_upstream AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --dma/read_master pcie_to_hibi_4x_sopc_burst_3/upstream arbiterlock, which is an e_assign
  dma_read_master_arbiterlock <= pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable AND dma_read_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_3_upstream_arb_share_counter_next_value);
  --dma/read_master pcie_to_hibi_4x_sopc_burst_3/upstream arbiterlock2, which is an e_assign
  dma_read_master_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable2 AND dma_read_master_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_any_continuerequest <= std_logic'('1');
  --dma_read_master_continuerequest continued request, which is an e_assign
  dma_read_master_continuerequest <= std_logic'('1');
  internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream AND NOT ((((NOT dma_read_master_read_n AND dma_read_master_chipselect)) AND ((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_read_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dma_read_master_latency_counter))))))) OR (dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register)))));
  --unique name for pcie_to_hibi_4x_sopc_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_move_on_to_next_transaction <= pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo;
  --the currently selected burstcount for pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 12);
  --burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream : burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_3_upstream_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_3_upstream_transaction_burst_count,
      empty => pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input14,
      clk => clk,
      data_in => pcie_to_hibi_4x_sopc_burst_3_upstream_selected_burstcount,
      read => pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input15,
      write => module_input16
    );

  module_input14 <= std_logic'('0');
  module_input15 <= std_logic'('0');
  module_input16 <= ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo) AND NOT ((pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount_fifo_empty));

  --pcie_to_hibi_4x_sopc_burst_3_upstream current burst minus one, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 12);
  --what to load in current_burst, for pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo))) = '1'), (pcie_to_hibi_4x_sopc_burst_3_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst) AND pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount_fifo_empty))) = '1'), (pcie_to_hibi_4x_sopc_burst_3_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst)) = '1'), (pcie_to_hibi_4x_sopc_burst_3_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst_minus_one))))), 12);
  --the current burst count for pcie_to_hibi_4x_sopc_burst_3_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa OR ((NOT pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo AND ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read)))))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst <= pcie_to_hibi_4x_sopc_burst_3_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read)) AND pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo) OR pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst)) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo <= p0_pcie_to_hibi_4x_sopc_burst_3_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(pcie_to_hibi_4x_sopc_burst_3_upstream_current_burst_minus_one)) AND pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream : rdv_fifo_for_dma_read_master_to_pcie_to_hibi_4x_sopc_burst_3_upstream_module
    port map(
      data_out => dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_3_upstream,
      empty => open,
      fifo_contains_ones_n => dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_3_upstream,
      full => open,
      clear_fifo => module_input17,
      clk => clk,
      data_in => internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream,
      read => pcie_to_hibi_4x_sopc_burst_3_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => dma_read_master_flush_qualified_exported,
      write => module_input18
    );

  module_input17 <= std_logic'('0');
  module_input18 <= in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read;

  dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register <= NOT dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --local readdatavalid dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_mux
  dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream <= ((pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid_from_sa AND dma_read_master_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_3_upstream)) AND NOT dma_read_master_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_3/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress <= dma_read_master_address_to_slave (15 DOWNTO 0);
  --master is always granted when requested
  internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --dma/read_master saved-grant pcie_to_hibi_4x_sopc_burst_3/upstream, which is an e_assign
  dma_read_master_saved_grant_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_3/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_3_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_3_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_3_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_3_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_3_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_3_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_3_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_3_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_3_upstream_write) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("0000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_3_upstream_read) AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 10);
  --pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_3_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_3_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_3_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_3_upstream_read <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --pcie_to_hibi_4x_sopc_burst_3_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_3_upstream_write <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_3_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(dma_read_master_address_to_slave,std_logic_vector'("00000000000000000000000000000011")) & A_ToStdLogicVector(dma_read_master_dbs_address(2)) & A_REP(std_logic'('0'), 2)), 14);
  --d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_read_cycle <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream AND ((NOT dma_read_master_read_n AND dma_read_master_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_3_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_3_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream)) = '1'), (std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --vhdl renameroo for output signals
  dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --vhdl renameroo for output signals
  dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream <= internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_3_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_3_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_3/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --dma/read_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream AND to_std_logic((((std_logic_vector'("000000000000000000000") & (dma_read_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("dma/read_master drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_3/upstream"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pcie_Control_Register_Access_end_xfer : IN STD_LOGIC;
                 signal pcie_Control_Register_Access_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Control_Register_Access_waitrequest_from_sa : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_last_time :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_is_granted_some_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access OR NOT pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access OR NOT pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access OR NOT ((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Control_Register_Access_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access OR NOT ((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_Control_Register_Access_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_3_downstream_address;
  --pcie_to_hibi_4x_sopc_burst_3_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_3_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcie_to_hibi_4x_sopc_burst_3_downstream_read_but_no_slave_selected <= (pcie_to_hibi_4x_sopc_burst_3_downstream_read AND pcie_to_hibi_4x_sopc_burst_3_downstream_run) AND NOT pcie_to_hibi_4x_sopc_burst_3_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_downstream_is_granted_some_slave <= pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid <= (pcie_to_hibi_4x_sopc_burst_3_downstream_read_but_no_slave_selected OR pre_flush_pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid) OR pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access;
  --pcie_to_hibi_4x_sopc_burst_3/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_3_downstream_readdata <= pcie_Control_Register_Access_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_3_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter <= p1_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pcie_to_hibi_4x_sopc_burst_3_downstream_run AND pcie_to_hibi_4x_sopc_burst_3_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_3_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_address_last_time <= std_logic_vector'("00000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_3_downstream_read OR pcie_to_hibi_4x_sopc_burst_3_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_3_downstream_address /= pcie_to_hibi_4x_sopc_burst_3_downstream_address_last_time))))) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_address did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount) /= std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable_last_time))))) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_read_last_time)))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_read did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_3_downstream_write_last_time)))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_write did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_3_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_3_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_3_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_3_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_3_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_3_downstream_write)) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("pcie_to_hibi_4x_sopc_burst_3_downstream_writedata did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module;


architecture europa of burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module;


architecture europa of rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcie_Rx_Interface_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_Rx_Interface_latency_counter : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal pcie_Rx_Interface_write : IN STD_LOGIC;
                 signal pcie_Rx_Interface_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_write : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator is
component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module;

component rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_4_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_upstream_write :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal p0_pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal pcie_Rx_Interface_arbiterlock :  STD_LOGIC;
                signal pcie_Rx_Interface_arbiterlock2 :  STD_LOGIC;
                signal pcie_Rx_Interface_continuerequest :  STD_LOGIC;
                signal pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_next_burst_count :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_selected_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pcie_to_hibi_4x_sopc_burst_4_upstream_from_pcie_Rx_Interface :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_pcie_to_hibi_4x_sopc_burst_4_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_4_upstream_readdata;
  internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream <= to_std_logic(((Std_Logic_Vector'(pcie_Rx_Interface_address_to_slave(31 DOWNTO 6) & std_logic_vector'("000000")) = std_logic_vector'("10000000000000000001000000000000")))) AND ((pcie_Rx_Interface_read OR pcie_Rx_Interface_write));
  --assign pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest;
  --assign pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((pcie_Rx_Interface_write)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 12);
  --pcie_to_hibi_4x_sopc_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_any_bursting_master_saved_grant <= pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_4_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 12);
  --pcie_to_hibi_4x_sopc_burst_4_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_4_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream <= pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_4_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream AND pcie_to_hibi_4x_sopc_burst_4_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_4_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_4_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_4_upstream AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie/Rx_Interface pcie_to_hibi_4x_sopc_burst_4/upstream arbiterlock, which is an e_assign
  pcie_Rx_Interface_arbiterlock <= pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable AND pcie_Rx_Interface_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_4_upstream_arb_share_counter_next_value);
  --pcie/Rx_Interface pcie_to_hibi_4x_sopc_burst_4/upstream arbiterlock2, which is an e_assign
  pcie_Rx_Interface_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable2 AND pcie_Rx_Interface_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_any_continuerequest <= std_logic'('1');
  --pcie_Rx_Interface_continuerequest continued request, which is an e_assign
  pcie_Rx_Interface_continuerequest <= std_logic'('1');
  internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream AND NOT ((pcie_Rx_Interface_read AND ((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_latency_counter))))))) OR (pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register)))));
  --unique name for pcie_to_hibi_4x_sopc_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_move_on_to_next_transaction <= pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo;
  --the currently selected burstcount for pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 10);
  --burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream : burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_4_upstream_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_4_upstream_transaction_burst_count,
      empty => pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input19,
      clk => clk,
      data_in => pcie_to_hibi_4x_sopc_burst_4_upstream_selected_burstcount,
      read => pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input20,
      write => module_input21
    );

  module_input19 <= std_logic'('0');
  module_input20 <= std_logic'('0');
  module_input21 <= ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo) AND NOT ((pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount_fifo_empty));

  --pcie_to_hibi_4x_sopc_burst_4_upstream current burst minus one, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 10);
  --what to load in current_burst, for pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo))) = '1'), pcie_to_hibi_4x_sopc_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst) AND pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount_fifo_empty))) = '1'), pcie_to_hibi_4x_sopc_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst)) = '1'), pcie_to_hibi_4x_sopc_burst_4_upstream_transaction_burst_count, pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst_minus_one)));
  --the current burst count for pcie_to_hibi_4x_sopc_burst_4_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst <= std_logic_vector'("0000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa OR ((NOT pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo AND ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read)))))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst <= pcie_to_hibi_4x_sopc_burst_4_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read)) AND pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo) OR pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst)) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo <= p0_pcie_to_hibi_4x_sopc_burst_4_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(pcie_to_hibi_4x_sopc_burst_4_upstream_current_burst_minus_one)) AND pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream : rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_4_upstream_module
    port map(
      data_out => pcie_Rx_Interface_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_4_upstream,
      empty => open,
      fifo_contains_ones_n => pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_4_upstream,
      full => open,
      clear_fifo => module_input22,
      clk => clk,
      data_in => internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream,
      read => pcie_to_hibi_4x_sopc_burst_4_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input23,
      write => module_input24
    );

  module_input22 <= std_logic'('0');
  module_input23 <= std_logic'('0');
  module_input24 <= in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read;

  pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register <= NOT pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --local readdatavalid pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_mux
  pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream <= pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid_from_sa;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_writedata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_writedata <= pcie_Rx_Interface_writedata (31 DOWNTO 0);
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_4/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress <= pcie_Rx_Interface_address_to_slave (6 DOWNTO 0);
  --master is always granted when requested
  internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --pcie/Rx_Interface saved-grant pcie_to_hibi_4x_sopc_burst_4/upstream, which is an e_assign
  pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_4/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_4_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_4_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_4_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_4_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_4_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_4_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_4_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_4_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_4_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_4_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 9);
  --pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter <= std_logic_vector'("000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_4_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_4_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_4_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_4_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_4_upstream_read <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream AND pcie_Rx_Interface_read;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_4_upstream_write <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream AND pcie_Rx_Interface_write;
  shifted_address_to_pcie_to_hibi_4x_sopc_burst_4_upstream_from_pcie_Rx_Interface <= pcie_Rx_Interface_address_to_slave;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_address <= A_EXT (A_SRL(shifted_address_to_pcie_to_hibi_4x_sopc_burst_4_upstream_from_pcie_Rx_Interface,std_logic_vector'("00000000000000000000000000000011")), 5);
  --d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_read_cycle <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream AND pcie_Rx_Interface_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_write_cycle <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream AND pcie_Rx_Interface_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_4_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_4_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream)) = '1'), (std_logic_vector'("000000000000000000000000") & (pcie_Rx_Interface_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 10);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_4_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_4_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_4/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie/Rx_Interface non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("pcie/Rx_Interface drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_4/upstream"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_dma_control_port_slave_end_xfer : IN STD_LOGIC;
                 signal dma_control_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_last_time :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave OR NOT pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave OR NOT ((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dma_control_port_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave OR NOT ((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dma_control_port_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_4_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave)))));
  --pcie_to_hibi_4x_sopc_burst_4/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_4_downstream_readdata <= dma_control_port_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_4_downstream_run;
  --latent max counter, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_4_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_address_last_time <= std_logic_vector'("00000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_4_downstream_read OR pcie_to_hibi_4x_sopc_burst_4_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_4_downstream_address /= pcie_to_hibi_4x_sopc_burst_4_downstream_address_last_time))))) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_address did not heed wait!!!"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount) /= std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable_last_time))))) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable did not heed wait!!!"));
          write(output, write_line63.all);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_read_last_time)))))) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_read did not heed wait!!!"));
          write(output, write_line64.all);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line65 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_4_downstream_write_last_time)))))) = '1' then 
          write(write_line65, now);
          write(write_line65, string'(": "));
          write(write_line65, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_write did not heed wait!!!"));
          write(output, write_line65.all);
          deallocate (write_line65);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_4_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_4_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_4_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line66 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_4_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_4_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_4_downstream_write)) = '1' then 
          write(write_line66, now);
          write(write_line66, string'(": "));
          write(write_line66, string'("pcie_to_hibi_4x_sopc_burst_4_downstream_writedata did not heed wait!!!"));
          write(output, write_line66.all);
          deallocate (write_line66);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module;


architecture europa of burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module;


architecture europa of rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcie_Rx_Interface_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pcie_Rx_Interface_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pcie_Rx_Interface_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_Rx_Interface_latency_counter : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read : IN STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal pcie_Rx_Interface_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : OUT STD_LOGIC;
                 signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_read : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_write : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator is
component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module;

component rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_5_upstream_read :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_upstream_write :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC;
                signal module_input29 :  STD_LOGIC;
                signal module_input30 :  STD_LOGIC;
                signal p0_pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal pcie_Rx_Interface_arbiterlock :  STD_LOGIC;
                signal pcie_Rx_Interface_arbiterlock2 :  STD_LOGIC;
                signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Rx_Interface_continuerequest :  STD_LOGIC;
                signal pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_allgrants :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_any_continuerequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_arb_counter_enable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_grant_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_read_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_write_cycle :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_master_qreq_vector :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_next_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_reg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_selected_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_write :  STD_LOGIC;
                signal wait_for_pcie_to_hibi_4x_sopc_burst_5_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer;
    end if;

  end process;

  pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream);
  --assign pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa = pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa <= pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid;
  --assign pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa = pcie_to_hibi_4x_sopc_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa <= pcie_to_hibi_4x_sopc_burst_5_upstream_readdata;
  internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream <= to_std_logic(((Std_Logic_Vector'(pcie_Rx_Interface_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND ((pcie_Rx_Interface_read OR pcie_Rx_Interface_write));
  --assign pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa = pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa <= pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter set values, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((pcie_Rx_Interface_write)) = '1'), (std_logic_vector'("0000000000000000000000") & (A_SLL(pcie_Rx_Interface_burstcount,std_logic_vector'("00000000000000000000000000000001")))), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 12);
  --pcie_to_hibi_4x_sopc_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_non_bursting_master_requests <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_any_bursting_master_saved_grant <= pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcie_to_hibi_4x_sopc_burst_5_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 12);
  --pcie_to_hibi_4x_sopc_burst_5_upstream_allgrants all slave grants, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_allgrants <= pcie_to_hibi_4x_sopc_burst_5_upstream_grant_vector;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer <= NOT ((pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read OR pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream <= pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer AND (((NOT pcie_to_hibi_4x_sopc_burst_5_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_to_hibi_4x_sopc_burst_5_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_non_bursting_master_requests));
  --pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_5_upstream_arb_counter_enable) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter <= pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pcie_to_hibi_4x_sopc_burst_5_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream)) OR ((end_xfer_arb_share_counter_term_pcie_to_hibi_4x_sopc_burst_5_upstream AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_non_bursting_master_requests)))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable <= or_reduce(pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcie/Rx_Interface pcie_to_hibi_4x_sopc_burst_5/upstream arbiterlock, which is an e_assign
  pcie_Rx_Interface_arbiterlock <= pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable AND pcie_Rx_Interface_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable2 <= or_reduce(pcie_to_hibi_4x_sopc_burst_5_upstream_arb_share_counter_next_value);
  --pcie/Rx_Interface pcie_to_hibi_4x_sopc_burst_5/upstream arbiterlock2, which is an e_assign
  pcie_Rx_Interface_arbiterlock2 <= pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable2 AND pcie_Rx_Interface_continuerequest;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_any_continuerequest <= std_logic'('1');
  --pcie_Rx_Interface_continuerequest continued request, which is an e_assign
  pcie_Rx_Interface_continuerequest <= std_logic'('1');
  internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream AND NOT ((pcie_Rx_Interface_read AND ((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_latency_counter))))))) OR (pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register)))));
  --unique name for pcie_to_hibi_4x_sopc_burst_5_upstream_move_on_to_next_transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_move_on_to_next_transaction <= pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo;
  --the currently selected burstcount for pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream : burstcount_fifo_for_pcie_to_hibi_4x_sopc_burst_5_upstream_module
    port map(
      data_out => pcie_to_hibi_4x_sopc_burst_5_upstream_transaction_burst_count,
      empty => pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input25,
      clk => clk,
      data_in => pcie_to_hibi_4x_sopc_burst_5_upstream_selected_burstcount,
      read => pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input26,
      write => module_input27
    );

  module_input25 <= std_logic'('0');
  module_input26 <= std_logic'('0');
  module_input27 <= ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo) AND NOT ((pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst AND pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount_fifo_empty));

  --pcie_to_hibi_4x_sopc_burst_5_upstream current burst minus one, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 11);
  --what to load in current_burst, for pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo))) = '1'), (pcie_to_hibi_4x_sopc_burst_5_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read) AND pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst) AND pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount_fifo_empty))) = '1'), (pcie_to_hibi_4x_sopc_burst_5_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst)) = '1'), (pcie_to_hibi_4x_sopc_burst_5_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst_minus_one))))), 11);
  --the current burst count for pcie_to_hibi_4x_sopc_burst_5_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa OR ((NOT pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo AND ((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read)))))) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst <= pcie_to_hibi_4x_sopc_burst_5_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read)) AND pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read)) AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo) OR pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst)) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo <= p0_pcie_to_hibi_4x_sopc_burst_5_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(pcie_to_hibi_4x_sopc_burst_5_upstream_current_burst_minus_one)) AND pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream : rdv_fifo_for_pcie_Rx_Interface_to_pcie_to_hibi_4x_sopc_burst_5_upstream_module
    port map(
      data_out => pcie_Rx_Interface_rdv_fifo_output_from_pcie_to_hibi_4x_sopc_burst_5_upstream,
      empty => open,
      fifo_contains_ones_n => pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_5_upstream,
      full => open,
      clear_fifo => module_input28,
      clk => clk,
      data_in => internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream,
      read => pcie_to_hibi_4x_sopc_burst_5_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input29,
      write => module_input30
    );

  module_input28 <= std_logic'('0');
  module_input29 <= std_logic'('0');
  module_input30 <= in_a_read_cycle AND NOT pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read;

  pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register <= NOT pcie_Rx_Interface_rdv_fifo_empty_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --local readdatavalid pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_mux
  pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream <= pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid_from_sa;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_writedata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_writedata <= pcie_Rx_Interface_dbs_write_32;
  --byteaddress mux for pcie_to_hibi_4x_sopc_burst_5/upstream, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress <= pcie_Rx_Interface_address_to_slave (26 DOWNTO 0);
  --master is always granted when requested
  internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --pcie/Rx_Interface saved-grant pcie_to_hibi_4x_sopc_burst_5/upstream, which is an e_assign
  pcie_Rx_Interface_saved_grant_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --allow new arb cycle for pcie_to_hibi_4x_sopc_burst_5/upstream, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pcie_to_hibi_4x_sopc_burst_5_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pcie_to_hibi_4x_sopc_burst_5_upstream_master_qreq_vector <= std_logic'('1');
  --pcie_to_hibi_4x_sopc_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer) = '1'), pcie_to_hibi_4x_sopc_burst_5_upstream_unreg_firsttransfer, pcie_to_hibi_4x_sopc_burst_5_upstream_reg_firsttransfer);
  --pcie_to_hibi_4x_sopc_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_unreg_firsttransfer <= NOT ((pcie_to_hibi_4x_sopc_burst_5_upstream_slavearbiterlockenable AND pcie_to_hibi_4x_sopc_burst_5_upstream_any_continuerequest));
  --pcie_to_hibi_4x_sopc_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_reg_firsttransfer <= pcie_to_hibi_4x_sopc_burst_5_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_5_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000") & (internal_pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_pcie_to_hibi_4x_sopc_burst_5_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 9);
  --pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter <= std_logic_vector'("000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer) = '1' then 
        pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter <= pcie_to_hibi_4x_sopc_burst_5_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_beginbursttransfer_internal <= pcie_to_hibi_4x_sopc_burst_5_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (pcie_to_hibi_4x_sopc_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --pcie_to_hibi_4x_sopc_burst_5_upstream_read assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_5_upstream_read <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_read;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_write assignment, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_5_upstream_write <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_write;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_address mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(pcie_Rx_Interface_address_to_slave,std_logic_vector'("00000000000000000000000000000011")) & A_ToStdLogicVector(pcie_Rx_Interface_dbs_address(2)) & A_REP(std_logic'('0'), 2)), 25);
  --d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer <= pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer;
    end if;

  end process;

  --pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_read <= pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_read_cycle AND internal_pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_read_cycle <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_read_cycle;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_waits_for_write <= pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_write_cycle AND internal_pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa;
  --pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_write_cycle <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream AND pcie_Rx_Interface_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcie_to_hibi_4x_sopc_burst_5_upstream_in_a_write_cycle;
  wait_for_pcie_to_hibi_4x_sopc_burst_5_upstream_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (internal_pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  (pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1(3), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1(2), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1(1), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1(0), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0(3), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0(2), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0(1), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0(0)) <= pcie_Rx_Interface_byteenable;
  internal_pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_dbs_address(2)))) = std_logic_vector'("00000000000000000000000000000000"))), pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_0, pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream_segment_1);
  --burstcount mux, which is an e_mux
  internal_pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 10);
  --debugaccess mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --vhdl renameroo for output signals
  pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream <= internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount <= internal_pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_upstream_read <= internal_pcie_to_hibi_4x_sopc_burst_5_upstream_read;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa <= internal_pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_upstream_write <= internal_pcie_to_hibi_4x_sopc_burst_5_upstream_write;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_5/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pcie/Rx_Interface non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line67 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (pcie_Rx_Interface_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line67, now);
          write(write_line67, string'(": "));
          write(write_line67, string'("pcie/Rx_Interface drove 0 on its 'burstcount' port while accessing slave pcie_to_hibi_4x_sopc_burst_5/upstream"));
          write(output, write_line67.all);
          deallocate (write_line67);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator is 
        port (
              -- inputs:
                 signal a2h_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal a2h_avalon_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal d1_a2h_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_read : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_write : IN STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n : OUT STD_LOGIC;
                 signal pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator;


architecture europa of pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_run :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_write_last_time :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave OR NOT pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave OR NOT ((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT a2h_avalon_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave OR NOT ((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT a2h_avalon_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave <= pcie_to_hibi_4x_sopc_burst_5_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave)))));
  --pcie_to_hibi_4x_sopc_burst_5/downstream readdata mux, which is an e_mux
  pcie_to_hibi_4x_sopc_burst_5_downstream_readdata <= a2h_avalon_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest <= NOT pcie_to_hibi_4x_sopc_burst_5_downstream_run;
  --latent max counter, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter <= std_logic'('0');
  --pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n assignment, which is an e_assign
  pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave;
  --vhdl renameroo for output signals
  pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest;
--synthesis translate_off
    --pcie_to_hibi_4x_sopc_burst_5_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_address_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_address;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest AND ((pcie_to_hibi_4x_sopc_burst_5_downstream_read OR pcie_to_hibi_4x_sopc_burst_5_downstream_write));
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line68 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_5_downstream_address /= pcie_to_hibi_4x_sopc_burst_5_downstream_address_last_time))))) = '1' then 
          write(write_line68, now);
          write(write_line68, string'(": "));
          write(write_line68, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_address did not heed wait!!!"));
          write(output, write_line68.all);
          deallocate (write_line68);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line69 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount) /= std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line69, now);
          write(write_line69, string'(": "));
          write(write_line69, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount did not heed wait!!!"));
          write(output, write_line69.all);
          deallocate (write_line69);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line70 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable /= pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable_last_time))))) = '1' then 
          write(write_line70, now);
          write(write_line70, string'(": "));
          write(write_line70, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable did not heed wait!!!"));
          write(output, write_line70.all);
          deallocate (write_line70);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_read_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_read;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line71 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_read) /= std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_read_last_time)))))) = '1' then 
          write(write_line71, now);
          write(write_line71, string'(": "));
          write(write_line71, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_read did not heed wait!!!"));
          write(output, write_line71.all);
          deallocate (write_line71);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_write_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_write;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line72 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_write) /= std_logic'(pcie_to_hibi_4x_sopc_burst_5_downstream_write_last_time)))))) = '1' then 
          write(write_line72, now);
          write(write_line72, string'(": "));
          write(write_line72, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_write did not heed wait!!!"));
          write(output, write_line72.all);
          deallocate (write_line72);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcie_to_hibi_4x_sopc_burst_5_downstream_writedata_last_time <= pcie_to_hibi_4x_sopc_burst_5_downstream_writedata;
      end if;

    end process;

    --pcie_to_hibi_4x_sopc_burst_5_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line73 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pcie_to_hibi_4x_sopc_burst_5_downstream_writedata /= pcie_to_hibi_4x_sopc_burst_5_downstream_writedata_last_time)))) AND pcie_to_hibi_4x_sopc_burst_5_downstream_write)) = '1' then 
          write(write_line73, now);
          write(write_line73, string'(": "));
          write(write_line73, string'("pcie_to_hibi_4x_sopc_burst_5_downstream_writedata did not heed wait!!!"));
          write(output, write_line73.all);
          deallocate (write_line73);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module;


architecture europa of pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pcie_to_hibi_4x_sopc is 
        port (
              -- 1) global signals:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_a2h
                 signal hibi_av_in_to_the_a2h : IN STD_LOGIC;
                 signal hibi_av_out_from_the_a2h : OUT STD_LOGIC;
                 signal hibi_comm_in_to_the_a2h : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal hibi_comm_out_from_the_a2h : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal hibi_data_in_to_the_a2h : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal hibi_data_out_from_the_a2h : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal hibi_empty_in_to_the_a2h : IN STD_LOGIC;
                 signal hibi_full_in_to_the_a2h : IN STD_LOGIC;
                 signal hibi_one_d_in_to_the_a2h : IN STD_LOGIC;
                 signal hibi_one_p_in_to_the_a2h : IN STD_LOGIC;
                 signal hibi_re_out_from_the_a2h : OUT STD_LOGIC;
                 signal hibi_we_out_from_the_a2h : OUT STD_LOGIC;

              -- the_pcie
                 signal clk125_out_pcie : OUT STD_LOGIC;
                 signal clk250_out_pcie : OUT STD_LOGIC;
                 signal clk500_out_pcie : OUT STD_LOGIC;
                 signal gxb_powerdown_pcie : IN STD_LOGIC;
                 signal pcie_rstn_pcie : IN STD_LOGIC;
                 signal phystatus_ext_pcie : IN STD_LOGIC;
                 signal pipe_mode_pcie : IN STD_LOGIC;
                 signal pll_powerdown_pcie : IN STD_LOGIC;
                 signal powerdown_ext_pcie : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal rate_ext_pcie : OUT STD_LOGIC;
                 signal reconfig_clk_pcie : IN STD_LOGIC;
                 signal reconfig_fromgxb_pcie : OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
                 signal reconfig_togxb_pcie : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal refclk_pcie : IN STD_LOGIC;
                 signal rx_in0_pcie : IN STD_LOGIC;
                 signal rx_in1_pcie : IN STD_LOGIC;
                 signal rx_in2_pcie : IN STD_LOGIC;
                 signal rx_in3_pcie : IN STD_LOGIC;
                 signal rxdata0_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rxdata1_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rxdata2_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rxdata3_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rxdatak0_ext_pcie : IN STD_LOGIC;
                 signal rxdatak1_ext_pcie : IN STD_LOGIC;
                 signal rxdatak2_ext_pcie : IN STD_LOGIC;
                 signal rxdatak3_ext_pcie : IN STD_LOGIC;
                 signal rxelecidle0_ext_pcie : IN STD_LOGIC;
                 signal rxelecidle1_ext_pcie : IN STD_LOGIC;
                 signal rxelecidle2_ext_pcie : IN STD_LOGIC;
                 signal rxelecidle3_ext_pcie : IN STD_LOGIC;
                 signal rxpolarity0_ext_pcie : OUT STD_LOGIC;
                 signal rxpolarity1_ext_pcie : OUT STD_LOGIC;
                 signal rxpolarity2_ext_pcie : OUT STD_LOGIC;
                 signal rxpolarity3_ext_pcie : OUT STD_LOGIC;
                 signal rxstatus0_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal rxstatus1_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal rxstatus2_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal rxstatus3_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal rxvalid0_ext_pcie : IN STD_LOGIC;
                 signal rxvalid1_ext_pcie : IN STD_LOGIC;
                 signal rxvalid2_ext_pcie : IN STD_LOGIC;
                 signal rxvalid3_ext_pcie : IN STD_LOGIC;
                 signal test_in_pcie : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal test_out_pcie : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal tx_out0_pcie : OUT STD_LOGIC;
                 signal tx_out1_pcie : OUT STD_LOGIC;
                 signal tx_out2_pcie : OUT STD_LOGIC;
                 signal tx_out3_pcie : OUT STD_LOGIC;
                 signal txcompl0_ext_pcie : OUT STD_LOGIC;
                 signal txcompl1_ext_pcie : OUT STD_LOGIC;
                 signal txcompl2_ext_pcie : OUT STD_LOGIC;
                 signal txcompl3_ext_pcie : OUT STD_LOGIC;
                 signal txdata0_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal txdata1_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal txdata2_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal txdata3_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal txdatak0_ext_pcie : OUT STD_LOGIC;
                 signal txdatak1_ext_pcie : OUT STD_LOGIC;
                 signal txdatak2_ext_pcie : OUT STD_LOGIC;
                 signal txdatak3_ext_pcie : OUT STD_LOGIC;
                 signal txdetectrx_ext_pcie : OUT STD_LOGIC;
                 signal txelecidle0_ext_pcie : OUT STD_LOGIC;
                 signal txelecidle1_ext_pcie : OUT STD_LOGIC;
                 signal txelecidle2_ext_pcie : OUT STD_LOGIC;
                 signal txelecidle3_ext_pcie : OUT STD_LOGIC
              );
end entity pcie_to_hibi_4x_sopc;


architecture europa of pcie_to_hibi_4x_sopc is
component a2h_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal a2h_avalon_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal a2h_avalon_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal a2h_avalon_slave_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal a2h_avalon_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal a2h_avalon_slave_read : OUT STD_LOGIC;
                    signal a2h_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal a2h_avalon_slave_reset_n : OUT STD_LOGIC;
                    signal a2h_avalon_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal a2h_avalon_slave_write : OUT STD_LOGIC;
                    signal a2h_avalon_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_a2h_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave : OUT STD_LOGIC
                 );
end component a2h_avalon_slave_arbitrator;

component a2h is 
           port (
                 -- inputs:
                    signal av_addr_in : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal av_byte_en_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal av_re_in : IN STD_LOGIC;
                    signal av_we_in : IN STD_LOGIC;
                    signal av_wr_data_in : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal hibi_av_in : IN STD_LOGIC;
                    signal hibi_comm_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal hibi_data_in : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal hibi_empty_in : IN STD_LOGIC;
                    signal hibi_full_in : IN STD_LOGIC;
                    signal hibi_one_d_in : IN STD_LOGIC;
                    signal hibi_one_p_in : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_rd_data_out : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_wait_req_out : OUT STD_LOGIC;
                    signal hibi_av_out : OUT STD_LOGIC;
                    signal hibi_comm_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal hibi_data_out : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal hibi_re_out : OUT STD_LOGIC;
                    signal hibi_we_out : OUT STD_LOGIC
                 );
end component a2h;

component dma_control_port_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_control_port_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_control_port_slave_readyfordata : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_dma_control_port_slave_end_xfer : OUT STD_LOGIC;
                    signal dma_control_port_slave_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_control_port_slave_chipselect : OUT STD_LOGIC;
                    signal dma_control_port_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_control_port_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal dma_control_port_slave_reset_n : OUT STD_LOGIC;
                    signal dma_control_port_slave_write_n : OUT STD_LOGIC;
                    signal dma_control_port_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave : OUT STD_LOGIC
                 );
end component dma_control_port_slave_arbitrator;

component dma_read_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer : IN STD_LOGIC;
                    signal dma_read_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_read_master_chipselect : IN STD_LOGIC;
                    signal dma_read_master_flush : IN STD_LOGIC;
                    signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                    signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                    signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                    signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal dma_read_master_read_n : IN STD_LOGIC;
                    signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream : IN STD_LOGIC;
                    signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal dma_read_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_read_master_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_read_master_flush_qualified_exported : OUT STD_LOGIC;
                    signal dma_read_master_latency_counter : OUT STD_LOGIC;
                    signal dma_read_master_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal dma_read_master_readdatavalid : OUT STD_LOGIC;
                    signal dma_read_master_waitrequest : OUT STD_LOGIC
                 );
end component dma_read_master_arbitrator;

component dma_write_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer : IN STD_LOGIC;
                    signal dma_write_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal dma_write_master_chipselect : IN STD_LOGIC;
                    signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                    signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                    signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                    signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                    signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream : IN STD_LOGIC;
                    signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream : IN STD_LOGIC;
                    signal dma_write_master_write_n : IN STD_LOGIC;
                    signal dma_write_master_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal dma_write_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_write_master_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_waitrequest : OUT STD_LOGIC
                 );
end component dma_write_master_arbitrator;

component dma is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_ctl_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_ctl_chipselect : IN STD_LOGIC;
                    signal dma_ctl_write_n : IN STD_LOGIC;
                    signal dma_ctl_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal read_endofpacket : IN STD_LOGIC;
                    signal read_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal read_readdatavalid : IN STD_LOGIC;
                    signal read_waitrequest : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;
                    signal write_endofpacket : IN STD_LOGIC;
                    signal write_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal dma_ctl_irq : OUT STD_LOGIC;
                    signal dma_ctl_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_ctl_readyfordata : OUT STD_LOGIC;
                    signal read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal read_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal read_chipselect : OUT STD_LOGIC;
                    signal read_flush : OUT STD_LOGIC;
                    signal read_read_n : OUT STD_LOGIC;
                    signal write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal write_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal write_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal write_chipselect : OUT STD_LOGIC;
                    signal write_write_n : OUT STD_LOGIC;
                    signal write_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
                 );
end component dma;

component pcie_Control_Register_Access_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcie_Control_Register_Access_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Control_Register_Access_waitrequest : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_Control_Register_Access_end_xfer : OUT STD_LOGIC;
                    signal pcie_Control_Register_Access_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal pcie_Control_Register_Access_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_Control_Register_Access_chipselect : OUT STD_LOGIC;
                    signal pcie_Control_Register_Access_read : OUT STD_LOGIC;
                    signal pcie_Control_Register_Access_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Control_Register_Access_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_Control_Register_Access_write : OUT STD_LOGIC;
                    signal pcie_Control_Register_Access_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access : OUT STD_LOGIC
                 );
end component pcie_Control_Register_Access_arbitrator;

component pcie_Tx_Interface_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcie_Tx_Interface_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_Tx_Interface_readdatavalid : IN STD_LOGIC;
                    signal pcie_Tx_Interface_waitrequest : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_Tx_Interface_end_xfer : OUT STD_LOGIC;
                    signal pcie_Tx_Interface_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal pcie_Tx_Interface_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_Tx_Interface_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_Tx_Interface_chipselect : OUT STD_LOGIC;
                    signal pcie_Tx_Interface_read : OUT STD_LOGIC;
                    signal pcie_Tx_Interface_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_Tx_Interface_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_Tx_Interface_write : OUT STD_LOGIC;
                    signal pcie_Tx_Interface_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface : OUT STD_LOGIC
                 );
end component pcie_Tx_Interface_arbitrator;

component pcie_Rx_Interface_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer : IN STD_LOGIC;
                    signal pcie_Rx_Interface_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream : IN STD_LOGIC;
                    signal pcie_Rx_Interface_write : IN STD_LOGIC;
                    signal pcie_Rx_Interface_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_Rx_Interface_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_dbs_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pcie_Rx_Interface_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_latency_counter : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_Rx_Interface_readdatavalid : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_reset_n : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_waitrequest : OUT STD_LOGIC
                 );
end component pcie_Rx_Interface_arbitrator;

component pcie is 
           port (
                 -- inputs:
                    signal AvlClk_i : IN STD_LOGIC;
                    signal CraAddress_i : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal CraByteEnable_i : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal CraChipSelect_i : IN STD_LOGIC;
                    signal CraRead : IN STD_LOGIC;
                    signal CraWrite : IN STD_LOGIC;
                    signal CraWriteData_i : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal RxmIrqNum_i : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal RxmIrq_i : IN STD_LOGIC;
                    signal RxmReadDataValid_i : IN STD_LOGIC;
                    signal RxmReadData_i : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal RxmWaitRequest_i : IN STD_LOGIC;
                    signal TxsAddress_i : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal TxsBurstCount_i : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal TxsByteEnable_i : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal TxsChipSelect_i : IN STD_LOGIC;
                    signal TxsRead_i : IN STD_LOGIC;
                    signal TxsWriteData_i : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal TxsWrite_i : IN STD_LOGIC;
                    signal cal_blk_clk : IN STD_LOGIC;
                    signal gxb_powerdown : IN STD_LOGIC;
                    signal pcie_rstn : IN STD_LOGIC;
                    signal phystatus_ext : IN STD_LOGIC;
                    signal pipe_mode : IN STD_LOGIC;
                    signal pll_powerdown : IN STD_LOGIC;
                    signal reconfig_clk : IN STD_LOGIC;
                    signal reconfig_togxb : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal refclk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal rx_in0 : IN STD_LOGIC;
                    signal rx_in1 : IN STD_LOGIC;
                    signal rx_in2 : IN STD_LOGIC;
                    signal rx_in3 : IN STD_LOGIC;
                    signal rxdata0_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata1_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata2_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata3_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdatak0_ext : IN STD_LOGIC;
                    signal rxdatak1_ext : IN STD_LOGIC;
                    signal rxdatak2_ext : IN STD_LOGIC;
                    signal rxdatak3_ext : IN STD_LOGIC;
                    signal rxelecidle0_ext : IN STD_LOGIC;
                    signal rxelecidle1_ext : IN STD_LOGIC;
                    signal rxelecidle2_ext : IN STD_LOGIC;
                    signal rxelecidle3_ext : IN STD_LOGIC;
                    signal rxstatus0_ext : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus1_ext : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus2_ext : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus3_ext : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxvalid0_ext : IN STD_LOGIC;
                    signal rxvalid1_ext : IN STD_LOGIC;
                    signal rxvalid2_ext : IN STD_LOGIC;
                    signal rxvalid3_ext : IN STD_LOGIC;
                    signal test_in : IN STD_LOGIC_VECTOR (39 DOWNTO 0);

                 -- outputs:
                    signal CraIrq_o : OUT STD_LOGIC;
                    signal CraReadData_o : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal CraWaitRequest_o : OUT STD_LOGIC;
                    signal RxmAddress_o : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal RxmBurstCount_o : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal RxmByteEnable_o : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal RxmRead_o : OUT STD_LOGIC;
                    signal RxmResetRequest_o : OUT STD_LOGIC;
                    signal RxmWriteData_o : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal RxmWrite_o : OUT STD_LOGIC;
                    signal TxsReadDataValid_o : OUT STD_LOGIC;
                    signal TxsReadData_o : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal TxsWaitRequest_o : OUT STD_LOGIC;
                    signal clk125_out : OUT STD_LOGIC;
                    signal clk250_out : OUT STD_LOGIC;
                    signal clk500_out : OUT STD_LOGIC;
                    signal powerdown_ext : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rate_ext : OUT STD_LOGIC;
                    signal reconfig_fromgxb : OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
                    signal rxpolarity0_ext : OUT STD_LOGIC;
                    signal rxpolarity1_ext : OUT STD_LOGIC;
                    signal rxpolarity2_ext : OUT STD_LOGIC;
                    signal rxpolarity3_ext : OUT STD_LOGIC;
                    signal test_out : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal tx_out0 : OUT STD_LOGIC;
                    signal tx_out1 : OUT STD_LOGIC;
                    signal tx_out2 : OUT STD_LOGIC;
                    signal tx_out3 : OUT STD_LOGIC;
                    signal txcompl0_ext : OUT STD_LOGIC;
                    signal txcompl1_ext : OUT STD_LOGIC;
                    signal txcompl2_ext : OUT STD_LOGIC;
                    signal txcompl3_ext : OUT STD_LOGIC;
                    signal txdata0_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata1_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata2_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata3_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdatak0_ext : OUT STD_LOGIC;
                    signal txdatak1_ext : OUT STD_LOGIC;
                    signal txdatak2_ext : OUT STD_LOGIC;
                    signal txdatak3_ext : OUT STD_LOGIC;
                    signal txdetectrx_ext : OUT STD_LOGIC;
                    signal txelecidle0_ext : OUT STD_LOGIC;
                    signal txelecidle1_ext : OUT STD_LOGIC;
                    signal txelecidle2_ext : OUT STD_LOGIC;
                    signal txelecidle3_ext : OUT STD_LOGIC
                 );
end component pcie;

component pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_read_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_read_master_chipselect : IN STD_LOGIC;
                    signal dma_read_master_flush_qualified_exported : IN STD_LOGIC;
                    signal dma_read_master_latency_counter : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal dma_read_master_read_n : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                    signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                    signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : OUT STD_LOGIC;
                    signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_upstream_write : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_Tx_Interface_end_xfer : IN STD_LOGIC;
                    signal pcie_Tx_Interface_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_Tx_Interface_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_address : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_0;

component pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_write_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal dma_write_master_chipselect : IN STD_LOGIC;
                    signal dma_write_master_write_n : IN STD_LOGIC;
                    signal dma_write_master_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                    signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                    signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                    signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_write : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_upstream_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
                 );
end component pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_Tx_Interface_end_xfer : IN STD_LOGIC;
                    signal pcie_Tx_Interface_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_Tx_Interface_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_address : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_1 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_1;

component pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_write_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_write_master_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal dma_write_master_chipselect : IN STD_LOGIC;
                    signal dma_write_master_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_write_master_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_write_master_write_n : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                    signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                    signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                    signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_write : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_Control_Register_Access_end_xfer : IN STD_LOGIC;
                    signal pcie_Control_Register_Access_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Control_Register_Access_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_2 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC;
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_2;

component pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dma_read_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dma_read_master_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal dma_read_master_chipselect : IN STD_LOGIC;
                    signal dma_read_master_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dma_read_master_flush_qualified_exported : IN STD_LOGIC;
                    signal dma_read_master_latency_counter : IN STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal dma_read_master_read_n : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                    signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                    signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                    signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register : OUT STD_LOGIC;
                    signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_upstream_write : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pcie_Control_Register_Access_end_xfer : IN STD_LOGIC;
                    signal pcie_Control_Register_Access_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Control_Register_Access_waitrequest_from_sa : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_3 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC;
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_3;

component pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcie_Rx_Interface_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_Rx_Interface_latency_counter : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal pcie_Rx_Interface_write : IN STD_LOGIC;
                    signal pcie_Rx_Interface_writedata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_write : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_dma_control_port_slave_end_xfer : IN STD_LOGIC;
                    signal dma_control_port_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_4 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC;
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_4;

component pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcie_Rx_Interface_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_Rx_Interface_byteenable : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pcie_Rx_Interface_dbs_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pcie_Rx_Interface_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_Rx_Interface_latency_counter : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read : IN STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal pcie_Rx_Interface_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register : OUT STD_LOGIC;
                    signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_read : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_write : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal a2h_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal a2h_avalon_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal d1_a2h_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_read : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_write : IN STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n : OUT STD_LOGIC;
                    signal pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator;

component pcie_to_hibi_4x_sopc_burst_5 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC;
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_burst_5;

component pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module;

                signal a2h_avalon_slave_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal a2h_avalon_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal a2h_avalon_slave_read :  STD_LOGIC;
                signal a2h_avalon_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal a2h_avalon_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal a2h_avalon_slave_reset_n :  STD_LOGIC;
                signal a2h_avalon_slave_waitrequest :  STD_LOGIC;
                signal a2h_avalon_slave_waitrequest_from_sa :  STD_LOGIC;
                signal a2h_avalon_slave_write :  STD_LOGIC;
                signal a2h_avalon_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clk_reset_n :  STD_LOGIC;
                signal d1_a2h_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_dma_control_port_slave_end_xfer :  STD_LOGIC;
                signal d1_pcie_Control_Register_Access_end_xfer :  STD_LOGIC;
                signal d1_pcie_Tx_Interface_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal dma_control_port_slave_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_control_port_slave_chipselect :  STD_LOGIC;
                signal dma_control_port_slave_irq :  STD_LOGIC;
                signal dma_control_port_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_control_port_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_control_port_slave_readyfordata :  STD_LOGIC;
                signal dma_control_port_slave_readyfordata_from_sa :  STD_LOGIC;
                signal dma_control_port_slave_reset_n :  STD_LOGIC;
                signal dma_control_port_slave_write_n :  STD_LOGIC;
                signal dma_control_port_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_read_master_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_read_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_read_master_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_read_master_chipselect :  STD_LOGIC;
                signal dma_read_master_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_read_master_endofpacket :  STD_LOGIC;
                signal dma_read_master_flush :  STD_LOGIC;
                signal dma_read_master_flush_qualified_exported :  STD_LOGIC;
                signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_latency_counter :  STD_LOGIC;
                signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register :  STD_LOGIC;
                signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register :  STD_LOGIC;
                signal dma_read_master_read_n :  STD_LOGIC;
                signal dma_read_master_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal dma_read_master_readdatavalid :  STD_LOGIC;
                signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream :  STD_LOGIC;
                signal dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream :  STD_LOGIC;
                signal dma_read_master_waitrequest :  STD_LOGIC;
                signal dma_write_master_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_write_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_write_master_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal dma_write_master_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal dma_write_master_chipselect :  STD_LOGIC;
                signal dma_write_master_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dma_write_master_dbs_write_32 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dma_write_master_endofpacket :  STD_LOGIC;
                signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream :  STD_LOGIC;
                signal dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream :  STD_LOGIC;
                signal dma_write_master_waitrequest :  STD_LOGIC;
                signal dma_write_master_write_n :  STD_LOGIC;
                signal dma_write_master_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal internal_clk125_out_pcie :  STD_LOGIC;
                signal internal_clk250_out_pcie :  STD_LOGIC;
                signal internal_clk500_out_pcie :  STD_LOGIC;
                signal internal_hibi_av_out_from_the_a2h :  STD_LOGIC;
                signal internal_hibi_comm_out_from_the_a2h :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_hibi_data_out_from_the_a2h :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_hibi_re_out_from_the_a2h :  STD_LOGIC;
                signal internal_hibi_we_out_from_the_a2h :  STD_LOGIC;
                signal internal_powerdown_ext_pcie :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_rate_ext_pcie :  STD_LOGIC;
                signal internal_reconfig_fromgxb_pcie :  STD_LOGIC_VECTOR (16 DOWNTO 0);
                signal internal_rxpolarity0_ext_pcie :  STD_LOGIC;
                signal internal_rxpolarity1_ext_pcie :  STD_LOGIC;
                signal internal_rxpolarity2_ext_pcie :  STD_LOGIC;
                signal internal_rxpolarity3_ext_pcie :  STD_LOGIC;
                signal internal_test_out_pcie :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal internal_tx_out0_pcie :  STD_LOGIC;
                signal internal_tx_out1_pcie :  STD_LOGIC;
                signal internal_tx_out2_pcie :  STD_LOGIC;
                signal internal_tx_out3_pcie :  STD_LOGIC;
                signal internal_txcompl0_ext_pcie :  STD_LOGIC;
                signal internal_txcompl1_ext_pcie :  STD_LOGIC;
                signal internal_txcompl2_ext_pcie :  STD_LOGIC;
                signal internal_txcompl3_ext_pcie :  STD_LOGIC;
                signal internal_txdata0_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_txdata1_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_txdata2_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_txdata3_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_txdatak0_ext_pcie :  STD_LOGIC;
                signal internal_txdatak1_ext_pcie :  STD_LOGIC;
                signal internal_txdatak2_ext_pcie :  STD_LOGIC;
                signal internal_txdatak3_ext_pcie :  STD_LOGIC;
                signal internal_txdetectrx_ext_pcie :  STD_LOGIC;
                signal internal_txelecidle0_ext_pcie :  STD_LOGIC;
                signal internal_txelecidle1_ext_pcie :  STD_LOGIC;
                signal internal_txelecidle2_ext_pcie :  STD_LOGIC;
                signal internal_txelecidle3_ext_pcie :  STD_LOGIC;
                signal module_input31 :  STD_LOGIC;
                signal pcie_Control_Register_Access_address :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_Control_Register_Access_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Control_Register_Access_chipselect :  STD_LOGIC;
                signal pcie_Control_Register_Access_irq :  STD_LOGIC;
                signal pcie_Control_Register_Access_read :  STD_LOGIC;
                signal pcie_Control_Register_Access_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Control_Register_Access_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Control_Register_Access_waitrequest :  STD_LOGIC;
                signal pcie_Control_Register_Access_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_Control_Register_Access_write :  STD_LOGIC;
                signal pcie_Control_Register_Access_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Rx_Interface_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Rx_Interface_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Rx_Interface_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Rx_Interface_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_Rx_Interface_dbs_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pcie_Rx_Interface_dbs_write_32 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_irq :  STD_LOGIC;
                signal pcie_Rx_Interface_irqnumber :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal pcie_Rx_Interface_latency_counter :  STD_LOGIC;
                signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_read :  STD_LOGIC;
                signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register :  STD_LOGIC;
                signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register :  STD_LOGIC;
                signal pcie_Rx_Interface_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_Rx_Interface_readdatavalid :  STD_LOGIC;
                signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream :  STD_LOGIC;
                signal pcie_Rx_Interface_reset_n :  STD_LOGIC;
                signal pcie_Rx_Interface_resetrequest :  STD_LOGIC;
                signal pcie_Rx_Interface_waitrequest :  STD_LOGIC;
                signal pcie_Rx_Interface_write :  STD_LOGIC;
                signal pcie_Rx_Interface_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_Tx_Interface_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal pcie_Tx_Interface_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_Tx_Interface_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_Tx_Interface_chipselect :  STD_LOGIC;
                signal pcie_Tx_Interface_read :  STD_LOGIC;
                signal pcie_Tx_Interface_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_Tx_Interface_readdata_from_sa :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_Tx_Interface_readdatavalid :  STD_LOGIC;
                signal pcie_Tx_Interface_waitrequest :  STD_LOGIC;
                signal pcie_Tx_Interface_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_Tx_Interface_write :  STD_LOGIC;
                signal pcie_Tx_Interface_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_4_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_read :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_write :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal reset_n_sources :  STD_LOGIC;

begin

  --the_a2h_avalon_slave, which is an e_instance
  the_a2h_avalon_slave : a2h_avalon_slave_arbitrator
    port map(
      a2h_avalon_slave_address => a2h_avalon_slave_address,
      a2h_avalon_slave_byteenable => a2h_avalon_slave_byteenable,
      a2h_avalon_slave_read => a2h_avalon_slave_read,
      a2h_avalon_slave_readdata_from_sa => a2h_avalon_slave_readdata_from_sa,
      a2h_avalon_slave_reset_n => a2h_avalon_slave_reset_n,
      a2h_avalon_slave_waitrequest_from_sa => a2h_avalon_slave_waitrequest_from_sa,
      a2h_avalon_slave_write => a2h_avalon_slave_write,
      a2h_avalon_slave_writedata => a2h_avalon_slave_writedata,
      d1_a2h_avalon_slave_end_xfer => d1_a2h_avalon_slave_end_xfer,
      pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave,
      a2h_avalon_slave_readdata => a2h_avalon_slave_readdata,
      a2h_avalon_slave_waitrequest => a2h_avalon_slave_waitrequest,
      clk => clk,
      pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_5_downstream_read => pcie_to_hibi_4x_sopc_burst_5_downstream_read,
      pcie_to_hibi_4x_sopc_burst_5_downstream_write => pcie_to_hibi_4x_sopc_burst_5_downstream_write,
      pcie_to_hibi_4x_sopc_burst_5_downstream_writedata => pcie_to_hibi_4x_sopc_burst_5_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_a2h, which is an e_ptf_instance
  the_a2h : a2h
    port map(
      av_rd_data_out => a2h_avalon_slave_readdata,
      av_wait_req_out => a2h_avalon_slave_waitrequest,
      hibi_av_out => internal_hibi_av_out_from_the_a2h,
      hibi_comm_out => internal_hibi_comm_out_from_the_a2h,
      hibi_data_out => internal_hibi_data_out_from_the_a2h,
      hibi_re_out => internal_hibi_re_out_from_the_a2h,
      hibi_we_out => internal_hibi_we_out_from_the_a2h,
      av_addr_in => a2h_avalon_slave_address,
      av_byte_en_in => a2h_avalon_slave_byteenable,
      av_re_in => a2h_avalon_slave_read,
      av_we_in => a2h_avalon_slave_write,
      av_wr_data_in => a2h_avalon_slave_writedata,
      clk => clk,
      hibi_av_in => hibi_av_in_to_the_a2h,
      hibi_comm_in => hibi_comm_in_to_the_a2h,
      hibi_data_in => hibi_data_in_to_the_a2h,
      hibi_empty_in => hibi_empty_in_to_the_a2h,
      hibi_full_in => hibi_full_in_to_the_a2h,
      hibi_one_d_in => hibi_one_d_in_to_the_a2h,
      hibi_one_p_in => hibi_one_p_in_to_the_a2h,
      rst_n => a2h_avalon_slave_reset_n
    );


  --the_dma_control_port_slave, which is an e_instance
  the_dma_control_port_slave : dma_control_port_slave_arbitrator
    port map(
      d1_dma_control_port_slave_end_xfer => d1_dma_control_port_slave_end_xfer,
      dma_control_port_slave_address => dma_control_port_slave_address,
      dma_control_port_slave_chipselect => dma_control_port_slave_chipselect,
      dma_control_port_slave_readdata_from_sa => dma_control_port_slave_readdata_from_sa,
      dma_control_port_slave_readyfordata_from_sa => dma_control_port_slave_readyfordata_from_sa,
      dma_control_port_slave_reset_n => dma_control_port_slave_reset_n,
      dma_control_port_slave_write_n => dma_control_port_slave_write_n,
      dma_control_port_slave_writedata => dma_control_port_slave_writedata,
      pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave,
      clk => clk,
      dma_control_port_slave_readdata => dma_control_port_slave_readdata,
      dma_control_port_slave_readyfordata => dma_control_port_slave_readyfordata,
      pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress,
      pcie_to_hibi_4x_sopc_burst_4_downstream_read => pcie_to_hibi_4x_sopc_burst_4_downstream_read,
      pcie_to_hibi_4x_sopc_burst_4_downstream_write => pcie_to_hibi_4x_sopc_burst_4_downstream_write,
      pcie_to_hibi_4x_sopc_burst_4_downstream_writedata => pcie_to_hibi_4x_sopc_burst_4_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_dma_read_master, which is an e_instance
  the_dma_read_master : dma_read_master_arbitrator
    port map(
      dma_read_master_address_to_slave => dma_read_master_address_to_slave,
      dma_read_master_dbs_address => dma_read_master_dbs_address,
      dma_read_master_flush_qualified_exported => dma_read_master_flush_qualified_exported,
      dma_read_master_latency_counter => dma_read_master_latency_counter,
      dma_read_master_readdata => dma_read_master_readdata,
      dma_read_master_readdatavalid => dma_read_master_readdatavalid,
      dma_read_master_waitrequest => dma_read_master_waitrequest,
      clk => clk,
      d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer,
      d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer,
      dma_read_master_address => dma_read_master_address,
      dma_read_master_burstcount => dma_read_master_burstcount,
      dma_read_master_chipselect => dma_read_master_chipselect,
      dma_read_master_flush => dma_read_master_flush,
      dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register,
      dma_read_master_read_n => dma_read_master_read_n,
      dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream,
      pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa,
      reset_n => clk_reset_n
    );


  --the_dma_write_master, which is an e_instance
  the_dma_write_master : dma_write_master_arbitrator
    port map(
      dma_write_master_address_to_slave => dma_write_master_address_to_slave,
      dma_write_master_dbs_address => dma_write_master_dbs_address,
      dma_write_master_dbs_write_32 => dma_write_master_dbs_write_32,
      dma_write_master_waitrequest => dma_write_master_waitrequest,
      clk => clk,
      d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer,
      d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer,
      dma_write_master_address => dma_write_master_address,
      dma_write_master_burstcount => dma_write_master_burstcount,
      dma_write_master_byteenable => dma_write_master_byteenable,
      dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_chipselect => dma_write_master_chipselect,
      dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream,
      dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream,
      dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream,
      dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_write_n => dma_write_master_write_n,
      dma_write_master_writedata => dma_write_master_writedata,
      pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa,
      reset_n => clk_reset_n
    );


  --the_dma, which is an e_ptf_instance
  the_dma : dma
    port map(
      dma_ctl_irq => dma_control_port_slave_irq,
      dma_ctl_readdata => dma_control_port_slave_readdata,
      dma_ctl_readyfordata => dma_control_port_slave_readyfordata,
      read_address => dma_read_master_address,
      read_burstcount => dma_read_master_burstcount,
      read_chipselect => dma_read_master_chipselect,
      read_flush => dma_read_master_flush,
      read_read_n => dma_read_master_read_n,
      write_address => dma_write_master_address,
      write_burstcount => dma_write_master_burstcount,
      write_byteenable => dma_write_master_byteenable,
      write_chipselect => dma_write_master_chipselect,
      write_write_n => dma_write_master_write_n,
      write_writedata => dma_write_master_writedata,
      clk => clk,
      dma_ctl_address => dma_control_port_slave_address,
      dma_ctl_chipselect => dma_control_port_slave_chipselect,
      dma_ctl_write_n => dma_control_port_slave_write_n,
      dma_ctl_writedata => dma_control_port_slave_writedata,
      read_endofpacket => dma_read_master_endofpacket,
      read_readdata => dma_read_master_readdata,
      read_readdatavalid => dma_read_master_readdatavalid,
      read_waitrequest => dma_read_master_waitrequest,
      system_reset_n => dma_control_port_slave_reset_n,
      write_endofpacket => dma_write_master_endofpacket,
      write_waitrequest => dma_write_master_waitrequest
    );


  --the_pcie_Control_Register_Access, which is an e_instance
  the_pcie_Control_Register_Access : pcie_Control_Register_Access_arbitrator
    port map(
      d1_pcie_Control_Register_Access_end_xfer => d1_pcie_Control_Register_Access_end_xfer,
      pcie_Control_Register_Access_address => pcie_Control_Register_Access_address,
      pcie_Control_Register_Access_byteenable => pcie_Control_Register_Access_byteenable,
      pcie_Control_Register_Access_chipselect => pcie_Control_Register_Access_chipselect,
      pcie_Control_Register_Access_read => pcie_Control_Register_Access_read,
      pcie_Control_Register_Access_readdata_from_sa => pcie_Control_Register_Access_readdata_from_sa,
      pcie_Control_Register_Access_waitrequest_from_sa => pcie_Control_Register_Access_waitrequest_from_sa,
      pcie_Control_Register_Access_write => pcie_Control_Register_Access_write,
      pcie_Control_Register_Access_writedata => pcie_Control_Register_Access_writedata,
      pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access,
      clk => clk,
      pcie_Control_Register_Access_readdata => pcie_Control_Register_Access_readdata,
      pcie_Control_Register_Access_waitrequest => pcie_Control_Register_Access_waitrequest,
      pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_2_downstream_read => pcie_to_hibi_4x_sopc_burst_2_downstream_read,
      pcie_to_hibi_4x_sopc_burst_2_downstream_write => pcie_to_hibi_4x_sopc_burst_2_downstream_write,
      pcie_to_hibi_4x_sopc_burst_2_downstream_writedata => pcie_to_hibi_4x_sopc_burst_2_downstream_writedata,
      pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_3_downstream_read => pcie_to_hibi_4x_sopc_burst_3_downstream_read,
      pcie_to_hibi_4x_sopc_burst_3_downstream_write => pcie_to_hibi_4x_sopc_burst_3_downstream_write,
      pcie_to_hibi_4x_sopc_burst_3_downstream_writedata => pcie_to_hibi_4x_sopc_burst_3_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_Tx_Interface, which is an e_instance
  the_pcie_Tx_Interface : pcie_Tx_Interface_arbitrator
    port map(
      d1_pcie_Tx_Interface_end_xfer => d1_pcie_Tx_Interface_end_xfer,
      pcie_Tx_Interface_address => pcie_Tx_Interface_address,
      pcie_Tx_Interface_burstcount => pcie_Tx_Interface_burstcount,
      pcie_Tx_Interface_byteenable => pcie_Tx_Interface_byteenable,
      pcie_Tx_Interface_chipselect => pcie_Tx_Interface_chipselect,
      pcie_Tx_Interface_read => pcie_Tx_Interface_read,
      pcie_Tx_Interface_readdata_from_sa => pcie_Tx_Interface_readdata_from_sa,
      pcie_Tx_Interface_waitrequest_from_sa => pcie_Tx_Interface_waitrequest_from_sa,
      pcie_Tx_Interface_write => pcie_Tx_Interface_write,
      pcie_Tx_Interface_writedata => pcie_Tx_Interface_writedata,
      pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register => pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register,
      pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register => pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register,
      pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface,
      clk => clk,
      pcie_Tx_Interface_readdata => pcie_Tx_Interface_readdata,
      pcie_Tx_Interface_readdatavalid => pcie_Tx_Interface_readdatavalid,
      pcie_Tx_Interface_waitrequest => pcie_Tx_Interface_waitrequest,
      pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read => pcie_to_hibi_4x_sopc_burst_0_downstream_read,
      pcie_to_hibi_4x_sopc_burst_0_downstream_write => pcie_to_hibi_4x_sopc_burst_0_downstream_write,
      pcie_to_hibi_4x_sopc_burst_0_downstream_writedata => pcie_to_hibi_4x_sopc_burst_0_downstream_writedata,
      pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare,
      pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read => pcie_to_hibi_4x_sopc_burst_1_downstream_read,
      pcie_to_hibi_4x_sopc_burst_1_downstream_write => pcie_to_hibi_4x_sopc_burst_1_downstream_write,
      pcie_to_hibi_4x_sopc_burst_1_downstream_writedata => pcie_to_hibi_4x_sopc_burst_1_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_Rx_Interface, which is an e_instance
  the_pcie_Rx_Interface : pcie_Rx_Interface_arbitrator
    port map(
      pcie_Rx_Interface_address_to_slave => pcie_Rx_Interface_address_to_slave,
      pcie_Rx_Interface_dbs_address => pcie_Rx_Interface_dbs_address,
      pcie_Rx_Interface_dbs_write_32 => pcie_Rx_Interface_dbs_write_32,
      pcie_Rx_Interface_latency_counter => pcie_Rx_Interface_latency_counter,
      pcie_Rx_Interface_readdata => pcie_Rx_Interface_readdata,
      pcie_Rx_Interface_readdatavalid => pcie_Rx_Interface_readdatavalid,
      pcie_Rx_Interface_reset_n => pcie_Rx_Interface_reset_n,
      pcie_Rx_Interface_waitrequest => pcie_Rx_Interface_waitrequest,
      clk => clk,
      d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer,
      d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer,
      pcie_Rx_Interface_address => pcie_Rx_Interface_address,
      pcie_Rx_Interface_burstcount => pcie_Rx_Interface_burstcount,
      pcie_Rx_Interface_byteenable => pcie_Rx_Interface_byteenable,
      pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_read => pcie_Rx_Interface_read,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register,
      pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_write => pcie_Rx_Interface_write,
      pcie_Rx_Interface_writedata => pcie_Rx_Interface_writedata,
      pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa,
      reset_n => clk_reset_n
    );


  --the_pcie, which is an e_ptf_instance
  the_pcie : pcie
    port map(
      CraIrq_o => pcie_Control_Register_Access_irq,
      CraReadData_o => pcie_Control_Register_Access_readdata,
      CraWaitRequest_o => pcie_Control_Register_Access_waitrequest,
      RxmAddress_o => pcie_Rx_Interface_address,
      RxmBurstCount_o => pcie_Rx_Interface_burstcount,
      RxmByteEnable_o => pcie_Rx_Interface_byteenable,
      RxmRead_o => pcie_Rx_Interface_read,
      RxmResetRequest_o => pcie_Rx_Interface_resetrequest,
      RxmWriteData_o => pcie_Rx_Interface_writedata,
      RxmWrite_o => pcie_Rx_Interface_write,
      TxsReadDataValid_o => pcie_Tx_Interface_readdatavalid,
      TxsReadData_o => pcie_Tx_Interface_readdata,
      TxsWaitRequest_o => pcie_Tx_Interface_waitrequest,
      clk125_out => internal_clk125_out_pcie,
      clk250_out => internal_clk250_out_pcie,
      clk500_out => internal_clk500_out_pcie,
      powerdown_ext => internal_powerdown_ext_pcie,
      rate_ext => internal_rate_ext_pcie,
      reconfig_fromgxb => internal_reconfig_fromgxb_pcie,
      rxpolarity0_ext => internal_rxpolarity0_ext_pcie,
      rxpolarity1_ext => internal_rxpolarity1_ext_pcie,
      rxpolarity2_ext => internal_rxpolarity2_ext_pcie,
      rxpolarity3_ext => internal_rxpolarity3_ext_pcie,
      test_out => internal_test_out_pcie,
      tx_out0 => internal_tx_out0_pcie,
      tx_out1 => internal_tx_out1_pcie,
      tx_out2 => internal_tx_out2_pcie,
      tx_out3 => internal_tx_out3_pcie,
      txcompl0_ext => internal_txcompl0_ext_pcie,
      txcompl1_ext => internal_txcompl1_ext_pcie,
      txcompl2_ext => internal_txcompl2_ext_pcie,
      txcompl3_ext => internal_txcompl3_ext_pcie,
      txdata0_ext => internal_txdata0_ext_pcie,
      txdata1_ext => internal_txdata1_ext_pcie,
      txdata2_ext => internal_txdata2_ext_pcie,
      txdata3_ext => internal_txdata3_ext_pcie,
      txdatak0_ext => internal_txdatak0_ext_pcie,
      txdatak1_ext => internal_txdatak1_ext_pcie,
      txdatak2_ext => internal_txdatak2_ext_pcie,
      txdatak3_ext => internal_txdatak3_ext_pcie,
      txdetectrx_ext => internal_txdetectrx_ext_pcie,
      txelecidle0_ext => internal_txelecidle0_ext_pcie,
      txelecidle1_ext => internal_txelecidle1_ext_pcie,
      txelecidle2_ext => internal_txelecidle2_ext_pcie,
      txelecidle3_ext => internal_txelecidle3_ext_pcie,
      AvlClk_i => clk,
      CraAddress_i => pcie_Control_Register_Access_address,
      CraByteEnable_i => pcie_Control_Register_Access_byteenable,
      CraChipSelect_i => pcie_Control_Register_Access_chipselect,
      CraRead => pcie_Control_Register_Access_read,
      CraWrite => pcie_Control_Register_Access_write,
      CraWriteData_i => pcie_Control_Register_Access_writedata,
      RxmIrqNum_i => pcie_Rx_Interface_irqnumber,
      RxmIrq_i => pcie_Rx_Interface_irq,
      RxmReadDataValid_i => pcie_Rx_Interface_readdatavalid,
      RxmReadData_i => pcie_Rx_Interface_readdata,
      RxmWaitRequest_i => pcie_Rx_Interface_waitrequest,
      TxsAddress_i => pcie_Tx_Interface_address,
      TxsBurstCount_i => pcie_Tx_Interface_burstcount,
      TxsByteEnable_i => pcie_Tx_Interface_byteenable,
      TxsChipSelect_i => pcie_Tx_Interface_chipselect,
      TxsRead_i => pcie_Tx_Interface_read,
      TxsWriteData_i => pcie_Tx_Interface_writedata,
      TxsWrite_i => pcie_Tx_Interface_write,
      cal_blk_clk => clk,
      gxb_powerdown => gxb_powerdown_pcie,
      pcie_rstn => pcie_rstn_pcie,
      phystatus_ext => phystatus_ext_pcie,
      pipe_mode => pipe_mode_pcie,
      pll_powerdown => pll_powerdown_pcie,
      reconfig_clk => reconfig_clk_pcie,
      reconfig_togxb => reconfig_togxb_pcie,
      refclk => refclk_pcie,
      reset_n => pcie_Rx_Interface_reset_n,
      rx_in0 => rx_in0_pcie,
      rx_in1 => rx_in1_pcie,
      rx_in2 => rx_in2_pcie,
      rx_in3 => rx_in3_pcie,
      rxdata0_ext => rxdata0_ext_pcie,
      rxdata1_ext => rxdata1_ext_pcie,
      rxdata2_ext => rxdata2_ext_pcie,
      rxdata3_ext => rxdata3_ext_pcie,
      rxdatak0_ext => rxdatak0_ext_pcie,
      rxdatak1_ext => rxdatak1_ext_pcie,
      rxdatak2_ext => rxdatak2_ext_pcie,
      rxdatak3_ext => rxdatak3_ext_pcie,
      rxelecidle0_ext => rxelecidle0_ext_pcie,
      rxelecidle1_ext => rxelecidle1_ext_pcie,
      rxelecidle2_ext => rxelecidle2_ext_pcie,
      rxelecidle3_ext => rxelecidle3_ext_pcie,
      rxstatus0_ext => rxstatus0_ext_pcie,
      rxstatus1_ext => rxstatus1_ext_pcie,
      rxstatus2_ext => rxstatus2_ext_pcie,
      rxstatus3_ext => rxstatus3_ext_pcie,
      rxvalid0_ext => rxvalid0_ext_pcie,
      rxvalid1_ext => rxvalid1_ext_pcie,
      rxvalid2_ext => rxvalid2_ext_pcie,
      rxvalid3_ext => rxvalid3_ext_pcie,
      test_in => test_in_pcie
    );


  --the_pcie_to_hibi_4x_sopc_burst_0_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_0_upstream : pcie_to_hibi_4x_sopc_burst_0_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_0_upstream_end_xfer,
      dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register,
      dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream => dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_0_upstream,
      pcie_to_hibi_4x_sopc_burst_0_upstream_address => pcie_to_hibi_4x_sopc_burst_0_upstream_address,
      pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_0_upstream_read => pcie_to_hibi_4x_sopc_burst_0_upstream_read,
      pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_0_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_0_upstream_write => pcie_to_hibi_4x_sopc_burst_0_upstream_write,
      clk => clk,
      dma_read_master_address_to_slave => dma_read_master_address_to_slave,
      dma_read_master_burstcount => dma_read_master_burstcount,
      dma_read_master_chipselect => dma_read_master_chipselect,
      dma_read_master_flush_qualified_exported => dma_read_master_flush_qualified_exported,
      dma_read_master_latency_counter => dma_read_master_latency_counter,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register,
      dma_read_master_read_n => dma_read_master_read_n,
      pcie_to_hibi_4x_sopc_burst_0_upstream_readdata => pcie_to_hibi_4x_sopc_burst_0_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_0_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_0_downstream : pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_0_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_0_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_0_downstream_readdata => pcie_to_hibi_4x_sopc_burst_0_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest,
      clk => clk,
      d1_pcie_Tx_Interface_end_xfer => d1_pcie_Tx_Interface_end_xfer,
      pcie_Tx_Interface_readdata_from_sa => pcie_Tx_Interface_readdata_from_sa,
      pcie_Tx_Interface_waitrequest_from_sa => pcie_Tx_Interface_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_0_downstream_address => pcie_to_hibi_4x_sopc_burst_0_downstream_address,
      pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_granted_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_qualified_request_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read => pcie_to_hibi_4x_sopc_burst_0_downstream_read,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register => pcie_to_hibi_4x_sopc_burst_0_downstream_read_data_valid_pcie_Tx_Interface_shift_register,
      pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_0_downstream_requests_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_0_downstream_write => pcie_to_hibi_4x_sopc_burst_0_downstream_write,
      pcie_to_hibi_4x_sopc_burst_0_downstream_writedata => pcie_to_hibi_4x_sopc_burst_0_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_0, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_0 : pcie_to_hibi_4x_sopc_burst_0
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_0_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_0_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_0_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_0_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_0_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_0_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_0_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_0_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_0_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_0_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_0_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_0_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_0_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_0_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_0_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_0_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_0_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_0_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_0_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_0_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_0_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_0_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_0_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_0_upstream_writedata
    );


  --the_pcie_to_hibi_4x_sopc_burst_1_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_1_upstream : pcie_to_hibi_4x_sopc_burst_1_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_1_upstream_end_xfer,
      dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_1_upstream,
      dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_1_upstream,
      dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream => dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_1_upstream,
      pcie_to_hibi_4x_sopc_burst_1_upstream_address => pcie_to_hibi_4x_sopc_burst_1_upstream_address,
      pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_1_upstream_read => pcie_to_hibi_4x_sopc_burst_1_upstream_read,
      pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa => pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa,
      pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_1_upstream_write => pcie_to_hibi_4x_sopc_burst_1_upstream_write,
      pcie_to_hibi_4x_sopc_burst_1_upstream_writedata => pcie_to_hibi_4x_sopc_burst_1_upstream_writedata,
      clk => clk,
      dma_write_master_address_to_slave => dma_write_master_address_to_slave,
      dma_write_master_burstcount => dma_write_master_burstcount,
      dma_write_master_byteenable => dma_write_master_byteenable,
      dma_write_master_chipselect => dma_write_master_chipselect,
      dma_write_master_write_n => dma_write_master_write_n,
      dma_write_master_writedata => dma_write_master_writedata,
      pcie_to_hibi_4x_sopc_burst_1_upstream_readdata => pcie_to_hibi_4x_sopc_burst_1_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_1_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_1_downstream : pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_1_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_1_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_1_downstream_readdata => pcie_to_hibi_4x_sopc_burst_1_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest,
      clk => clk,
      d1_pcie_Tx_Interface_end_xfer => d1_pcie_Tx_Interface_end_xfer,
      pcie_Tx_Interface_readdata_from_sa => pcie_Tx_Interface_readdata_from_sa,
      pcie_Tx_Interface_waitrequest_from_sa => pcie_Tx_Interface_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_1_downstream_address => pcie_to_hibi_4x_sopc_burst_1_downstream_address,
      pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_granted_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_qualified_request_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read => pcie_to_hibi_4x_sopc_burst_1_downstream_read,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register => pcie_to_hibi_4x_sopc_burst_1_downstream_read_data_valid_pcie_Tx_Interface_shift_register,
      pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface => pcie_to_hibi_4x_sopc_burst_1_downstream_requests_pcie_Tx_Interface,
      pcie_to_hibi_4x_sopc_burst_1_downstream_write => pcie_to_hibi_4x_sopc_burst_1_downstream_write,
      pcie_to_hibi_4x_sopc_burst_1_downstream_writedata => pcie_to_hibi_4x_sopc_burst_1_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_1, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_1 : pcie_to_hibi_4x_sopc_burst_1
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_1_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_1_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_1_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_1_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_1_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_1_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_1_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_1_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_1_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_1_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_1_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_1_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_1_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_1_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_1_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_1_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_1_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_1_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_1_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_1_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_1_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_1_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_1_upstream_writedata
    );


  --the_pcie_to_hibi_4x_sopc_burst_2_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_2_upstream : pcie_to_hibi_4x_sopc_burst_2_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_2_upstream_end_xfer,
      dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_byteenable_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_granted_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_qualified_request_pcie_to_hibi_4x_sopc_burst_2_upstream,
      dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream => dma_write_master_requests_pcie_to_hibi_4x_sopc_burst_2_upstream,
      pcie_to_hibi_4x_sopc_burst_2_upstream_address => pcie_to_hibi_4x_sopc_burst_2_upstream_address,
      pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_2_upstream_read => pcie_to_hibi_4x_sopc_burst_2_upstream_read,
      pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa => pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa,
      pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_2_upstream_write => pcie_to_hibi_4x_sopc_burst_2_upstream_write,
      pcie_to_hibi_4x_sopc_burst_2_upstream_writedata => pcie_to_hibi_4x_sopc_burst_2_upstream_writedata,
      clk => clk,
      dma_write_master_address_to_slave => dma_write_master_address_to_slave,
      dma_write_master_burstcount => dma_write_master_burstcount,
      dma_write_master_byteenable => dma_write_master_byteenable,
      dma_write_master_chipselect => dma_write_master_chipselect,
      dma_write_master_dbs_address => dma_write_master_dbs_address,
      dma_write_master_dbs_write_32 => dma_write_master_dbs_write_32,
      dma_write_master_write_n => dma_write_master_write_n,
      pcie_to_hibi_4x_sopc_burst_2_upstream_readdata => pcie_to_hibi_4x_sopc_burst_2_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_2_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_2_downstream : pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_2_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_2_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_2_downstream_readdata => pcie_to_hibi_4x_sopc_burst_2_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest,
      clk => clk,
      d1_pcie_Control_Register_Access_end_xfer => d1_pcie_Control_Register_Access_end_xfer,
      pcie_Control_Register_Access_readdata_from_sa => pcie_Control_Register_Access_readdata_from_sa,
      pcie_Control_Register_Access_waitrequest_from_sa => pcie_Control_Register_Access_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_2_downstream_address => pcie_to_hibi_4x_sopc_burst_2_downstream_address,
      pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_granted_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_qualified_request_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_read => pcie_to_hibi_4x_sopc_burst_2_downstream_read,
      pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_read_data_valid_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_2_downstream_requests_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_2_downstream_write => pcie_to_hibi_4x_sopc_burst_2_downstream_write,
      pcie_to_hibi_4x_sopc_burst_2_downstream_writedata => pcie_to_hibi_4x_sopc_burst_2_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_2, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_2 : pcie_to_hibi_4x_sopc_burst_2
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_2_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_2_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_2_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_2_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_2_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_2_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_2_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_2_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_2_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_2_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_2_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_2_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_2_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_2_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_2_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_2_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_2_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_2_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_2_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_2_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_2_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_2_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_2_upstream_writedata
    );


  --the_pcie_to_hibi_4x_sopc_burst_3_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_3_upstream : pcie_to_hibi_4x_sopc_burst_3_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_3_upstream_end_xfer,
      dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_granted_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_qualified_request_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_3_upstream_shift_register,
      dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream => dma_read_master_requests_pcie_to_hibi_4x_sopc_burst_3_upstream,
      pcie_to_hibi_4x_sopc_burst_3_upstream_address => pcie_to_hibi_4x_sopc_burst_3_upstream_address,
      pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_3_upstream_read => pcie_to_hibi_4x_sopc_burst_3_upstream_read,
      pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_3_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_3_upstream_write => pcie_to_hibi_4x_sopc_burst_3_upstream_write,
      clk => clk,
      dma_read_master_address_to_slave => dma_read_master_address_to_slave,
      dma_read_master_burstcount => dma_read_master_burstcount,
      dma_read_master_chipselect => dma_read_master_chipselect,
      dma_read_master_dbs_address => dma_read_master_dbs_address,
      dma_read_master_flush_qualified_exported => dma_read_master_flush_qualified_exported,
      dma_read_master_latency_counter => dma_read_master_latency_counter,
      dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register => dma_read_master_read_data_valid_pcie_to_hibi_4x_sopc_burst_0_upstream_shift_register,
      dma_read_master_read_n => dma_read_master_read_n,
      pcie_to_hibi_4x_sopc_burst_3_upstream_readdata => pcie_to_hibi_4x_sopc_burst_3_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_3_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_3_downstream : pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_3_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_3_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_3_downstream_readdata => pcie_to_hibi_4x_sopc_burst_3_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest,
      clk => clk,
      d1_pcie_Control_Register_Access_end_xfer => d1_pcie_Control_Register_Access_end_xfer,
      pcie_Control_Register_Access_readdata_from_sa => pcie_Control_Register_Access_readdata_from_sa,
      pcie_Control_Register_Access_waitrequest_from_sa => pcie_Control_Register_Access_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_3_downstream_address => pcie_to_hibi_4x_sopc_burst_3_downstream_address,
      pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_granted_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_qualified_request_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_read => pcie_to_hibi_4x_sopc_burst_3_downstream_read,
      pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_read_data_valid_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access => pcie_to_hibi_4x_sopc_burst_3_downstream_requests_pcie_Control_Register_Access,
      pcie_to_hibi_4x_sopc_burst_3_downstream_write => pcie_to_hibi_4x_sopc_burst_3_downstream_write,
      pcie_to_hibi_4x_sopc_burst_3_downstream_writedata => pcie_to_hibi_4x_sopc_burst_3_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_3, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_3 : pcie_to_hibi_4x_sopc_burst_3
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_3_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_3_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_3_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_3_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_3_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_3_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_3_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_3_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_3_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_3_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_3_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_3_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_3_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_3_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_3_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_3_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_3_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_3_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_3_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_3_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_3_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_3_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_3_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_3_upstream_writedata
    );


  --the_pcie_to_hibi_4x_sopc_burst_4_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_4_upstream : pcie_to_hibi_4x_sopc_burst_4_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_4_upstream_end_xfer,
      pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register,
      pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream => pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_4_upstream,
      pcie_to_hibi_4x_sopc_burst_4_upstream_address => pcie_to_hibi_4x_sopc_burst_4_upstream_address,
      pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_4_upstream_read => pcie_to_hibi_4x_sopc_burst_4_upstream_read,
      pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_4_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_4_upstream_write => pcie_to_hibi_4x_sopc_burst_4_upstream_write,
      pcie_to_hibi_4x_sopc_burst_4_upstream_writedata => pcie_to_hibi_4x_sopc_burst_4_upstream_writedata,
      clk => clk,
      pcie_Rx_Interface_address_to_slave => pcie_Rx_Interface_address_to_slave,
      pcie_Rx_Interface_burstcount => pcie_Rx_Interface_burstcount,
      pcie_Rx_Interface_byteenable => pcie_Rx_Interface_byteenable,
      pcie_Rx_Interface_latency_counter => pcie_Rx_Interface_latency_counter,
      pcie_Rx_Interface_read => pcie_Rx_Interface_read,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register,
      pcie_Rx_Interface_write => pcie_Rx_Interface_write,
      pcie_Rx_Interface_writedata => pcie_Rx_Interface_writedata,
      pcie_to_hibi_4x_sopc_burst_4_upstream_readdata => pcie_to_hibi_4x_sopc_burst_4_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_4_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_4_downstream : pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_4_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_4_downstream_readdata => pcie_to_hibi_4x_sopc_burst_4_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest,
      clk => clk,
      d1_dma_control_port_slave_end_xfer => d1_dma_control_port_slave_end_xfer,
      dma_control_port_slave_readdata_from_sa => dma_control_port_slave_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_4_downstream_address => pcie_to_hibi_4x_sopc_burst_4_downstream_address,
      pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_granted_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_qualified_request_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_read => pcie_to_hibi_4x_sopc_burst_4_downstream_read,
      pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_read_data_valid_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave => pcie_to_hibi_4x_sopc_burst_4_downstream_requests_dma_control_port_slave,
      pcie_to_hibi_4x_sopc_burst_4_downstream_write => pcie_to_hibi_4x_sopc_burst_4_downstream_write,
      pcie_to_hibi_4x_sopc_burst_4_downstream_writedata => pcie_to_hibi_4x_sopc_burst_4_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_4, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_4 : pcie_to_hibi_4x_sopc_burst_4
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_4_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_4_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_4_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_4_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_4_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_4_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_4_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_4_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_4_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_4_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_4_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_4_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_4_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_4_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_4_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_4_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_4_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_4_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_4_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_4_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_4_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_4_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_4_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_4_upstream_writedata
    );


  --the_pcie_to_hibi_4x_sopc_burst_5_upstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_5_upstream : pcie_to_hibi_4x_sopc_burst_5_upstream_arbitrator
    port map(
      d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer => d1_pcie_to_hibi_4x_sopc_burst_5_upstream_end_xfer,
      pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_byteenable_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_granted_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_qualified_request_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_5_upstream_shift_register,
      pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream => pcie_Rx_Interface_requests_pcie_to_hibi_4x_sopc_burst_5_upstream,
      pcie_to_hibi_4x_sopc_burst_5_upstream_address => pcie_to_hibi_4x_sopc_burst_5_upstream_address,
      pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount => pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress => pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress,
      pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable => pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess,
      pcie_to_hibi_4x_sopc_burst_5_upstream_read => pcie_to_hibi_4x_sopc_burst_5_upstream_read,
      pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa => pcie_to_hibi_4x_sopc_burst_5_upstream_readdata_from_sa,
      pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa => pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest_from_sa,
      pcie_to_hibi_4x_sopc_burst_5_upstream_write => pcie_to_hibi_4x_sopc_burst_5_upstream_write,
      pcie_to_hibi_4x_sopc_burst_5_upstream_writedata => pcie_to_hibi_4x_sopc_burst_5_upstream_writedata,
      clk => clk,
      pcie_Rx_Interface_address_to_slave => pcie_Rx_Interface_address_to_slave,
      pcie_Rx_Interface_burstcount => pcie_Rx_Interface_burstcount,
      pcie_Rx_Interface_byteenable => pcie_Rx_Interface_byteenable,
      pcie_Rx_Interface_dbs_address => pcie_Rx_Interface_dbs_address,
      pcie_Rx_Interface_dbs_write_32 => pcie_Rx_Interface_dbs_write_32,
      pcie_Rx_Interface_latency_counter => pcie_Rx_Interface_latency_counter,
      pcie_Rx_Interface_read => pcie_Rx_Interface_read,
      pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register => pcie_Rx_Interface_read_data_valid_pcie_to_hibi_4x_sopc_burst_4_upstream_shift_register,
      pcie_Rx_Interface_write => pcie_Rx_Interface_write,
      pcie_to_hibi_4x_sopc_burst_5_upstream_readdata => pcie_to_hibi_4x_sopc_burst_5_upstream_readdata,
      pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_5_downstream, which is an e_instance
  the_pcie_to_hibi_4x_sopc_burst_5_downstream : pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrator
    port map(
      pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_address_to_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter => pcie_to_hibi_4x_sopc_burst_5_downstream_latency_counter,
      pcie_to_hibi_4x_sopc_burst_5_downstream_readdata => pcie_to_hibi_4x_sopc_burst_5_downstream_readdata,
      pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid,
      pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n => pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n,
      pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest,
      a2h_avalon_slave_readdata_from_sa => a2h_avalon_slave_readdata_from_sa,
      a2h_avalon_slave_waitrequest_from_sa => a2h_avalon_slave_waitrequest_from_sa,
      clk => clk,
      d1_a2h_avalon_slave_end_xfer => d1_a2h_avalon_slave_end_xfer,
      pcie_to_hibi_4x_sopc_burst_5_downstream_address => pcie_to_hibi_4x_sopc_burst_5_downstream_address,
      pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount => pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount,
      pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable => pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable,
      pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_granted_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_qualified_request_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_read => pcie_to_hibi_4x_sopc_burst_5_downstream_read,
      pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_read_data_valid_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave => pcie_to_hibi_4x_sopc_burst_5_downstream_requests_a2h_avalon_slave,
      pcie_to_hibi_4x_sopc_burst_5_downstream_write => pcie_to_hibi_4x_sopc_burst_5_downstream_write,
      pcie_to_hibi_4x_sopc_burst_5_downstream_writedata => pcie_to_hibi_4x_sopc_burst_5_downstream_writedata,
      reset_n => clk_reset_n
    );


  --the_pcie_to_hibi_4x_sopc_burst_5, which is an e_ptf_instance
  the_pcie_to_hibi_4x_sopc_burst_5 : pcie_to_hibi_4x_sopc_burst_5
    port map(
      downstream_address => pcie_to_hibi_4x_sopc_burst_5_downstream_address,
      downstream_arbitrationshare => pcie_to_hibi_4x_sopc_burst_5_downstream_arbitrationshare,
      downstream_burstcount => pcie_to_hibi_4x_sopc_burst_5_downstream_burstcount,
      downstream_byteenable => pcie_to_hibi_4x_sopc_burst_5_downstream_byteenable,
      downstream_debugaccess => pcie_to_hibi_4x_sopc_burst_5_downstream_debugaccess,
      downstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_5_downstream_nativeaddress,
      downstream_read => pcie_to_hibi_4x_sopc_burst_5_downstream_read,
      downstream_write => pcie_to_hibi_4x_sopc_burst_5_downstream_write,
      downstream_writedata => pcie_to_hibi_4x_sopc_burst_5_downstream_writedata,
      upstream_readdata => pcie_to_hibi_4x_sopc_burst_5_upstream_readdata,
      upstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_5_upstream_readdatavalid,
      upstream_waitrequest => pcie_to_hibi_4x_sopc_burst_5_upstream_waitrequest,
      clk => clk,
      downstream_readdata => pcie_to_hibi_4x_sopc_burst_5_downstream_readdata,
      downstream_readdatavalid => pcie_to_hibi_4x_sopc_burst_5_downstream_readdatavalid,
      downstream_waitrequest => pcie_to_hibi_4x_sopc_burst_5_downstream_waitrequest,
      reset_n => pcie_to_hibi_4x_sopc_burst_5_downstream_reset_n,
      upstream_address => pcie_to_hibi_4x_sopc_burst_5_upstream_byteaddress,
      upstream_burstcount => pcie_to_hibi_4x_sopc_burst_5_upstream_burstcount,
      upstream_byteenable => pcie_to_hibi_4x_sopc_burst_5_upstream_byteenable,
      upstream_debugaccess => pcie_to_hibi_4x_sopc_burst_5_upstream_debugaccess,
      upstream_nativeaddress => pcie_to_hibi_4x_sopc_burst_5_upstream_address,
      upstream_read => pcie_to_hibi_4x_sopc_burst_5_upstream_read,
      upstream_write => pcie_to_hibi_4x_sopc_burst_5_upstream_write,
      upstream_writedata => pcie_to_hibi_4x_sopc_burst_5_upstream_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  pcie_to_hibi_4x_sopc_reset_clk_domain_synch : pcie_to_hibi_4x_sopc_reset_clk_domain_synch_module
    port map(
      data_out => clk_reset_n,
      clk => clk,
      data_in => module_input31,
      reset_n => reset_n_sources
    );

  module_input31 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_resetrequest)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_resetrequest)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_resetrequest)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcie_Rx_Interface_resetrequest))))));
  --dma_read_master_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  dma_read_master_endofpacket <= std_logic'('0');
  --dma_write_master_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  dma_write_master_endofpacket <= std_logic'('0');
  --pcie_Rx_Interface_irq of type irq does not connect to anything so wire it to default (0)
  pcie_Rx_Interface_irq <= std_logic'('0');
  --pcie_Rx_Interface_irqnumber of type irqnumber does not connect to anything so wire it to default (0)
  pcie_Rx_Interface_irqnumber <= std_logic_vector'("000000");
  --pcie_to_hibi_4x_sopc_burst_0_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  pcie_to_hibi_4x_sopc_burst_0_upstream_writedata <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000");
  --pcie_to_hibi_4x_sopc_burst_3_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  pcie_to_hibi_4x_sopc_burst_3_upstream_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --vhdl renameroo for output signals
  clk125_out_pcie <= internal_clk125_out_pcie;
  --vhdl renameroo for output signals
  clk250_out_pcie <= internal_clk250_out_pcie;
  --vhdl renameroo for output signals
  clk500_out_pcie <= internal_clk500_out_pcie;
  --vhdl renameroo for output signals
  hibi_av_out_from_the_a2h <= internal_hibi_av_out_from_the_a2h;
  --vhdl renameroo for output signals
  hibi_comm_out_from_the_a2h <= internal_hibi_comm_out_from_the_a2h;
  --vhdl renameroo for output signals
  hibi_data_out_from_the_a2h <= internal_hibi_data_out_from_the_a2h;
  --vhdl renameroo for output signals
  hibi_re_out_from_the_a2h <= internal_hibi_re_out_from_the_a2h;
  --vhdl renameroo for output signals
  hibi_we_out_from_the_a2h <= internal_hibi_we_out_from_the_a2h;
  --vhdl renameroo for output signals
  powerdown_ext_pcie <= internal_powerdown_ext_pcie;
  --vhdl renameroo for output signals
  rate_ext_pcie <= internal_rate_ext_pcie;
  --vhdl renameroo for output signals
  reconfig_fromgxb_pcie <= internal_reconfig_fromgxb_pcie;
  --vhdl renameroo for output signals
  rxpolarity0_ext_pcie <= internal_rxpolarity0_ext_pcie;
  --vhdl renameroo for output signals
  rxpolarity1_ext_pcie <= internal_rxpolarity1_ext_pcie;
  --vhdl renameroo for output signals
  rxpolarity2_ext_pcie <= internal_rxpolarity2_ext_pcie;
  --vhdl renameroo for output signals
  rxpolarity3_ext_pcie <= internal_rxpolarity3_ext_pcie;
  --vhdl renameroo for output signals
  test_out_pcie <= internal_test_out_pcie;
  --vhdl renameroo for output signals
  tx_out0_pcie <= internal_tx_out0_pcie;
  --vhdl renameroo for output signals
  tx_out1_pcie <= internal_tx_out1_pcie;
  --vhdl renameroo for output signals
  tx_out2_pcie <= internal_tx_out2_pcie;
  --vhdl renameroo for output signals
  tx_out3_pcie <= internal_tx_out3_pcie;
  --vhdl renameroo for output signals
  txcompl0_ext_pcie <= internal_txcompl0_ext_pcie;
  --vhdl renameroo for output signals
  txcompl1_ext_pcie <= internal_txcompl1_ext_pcie;
  --vhdl renameroo for output signals
  txcompl2_ext_pcie <= internal_txcompl2_ext_pcie;
  --vhdl renameroo for output signals
  txcompl3_ext_pcie <= internal_txcompl3_ext_pcie;
  --vhdl renameroo for output signals
  txdata0_ext_pcie <= internal_txdata0_ext_pcie;
  --vhdl renameroo for output signals
  txdata1_ext_pcie <= internal_txdata1_ext_pcie;
  --vhdl renameroo for output signals
  txdata2_ext_pcie <= internal_txdata2_ext_pcie;
  --vhdl renameroo for output signals
  txdata3_ext_pcie <= internal_txdata3_ext_pcie;
  --vhdl renameroo for output signals
  txdatak0_ext_pcie <= internal_txdatak0_ext_pcie;
  --vhdl renameroo for output signals
  txdatak1_ext_pcie <= internal_txdatak1_ext_pcie;
  --vhdl renameroo for output signals
  txdatak2_ext_pcie <= internal_txdatak2_ext_pcie;
  --vhdl renameroo for output signals
  txdatak3_ext_pcie <= internal_txdatak3_ext_pcie;
  --vhdl renameroo for output signals
  txdetectrx_ext_pcie <= internal_txdetectrx_ext_pcie;
  --vhdl renameroo for output signals
  txelecidle0_ext_pcie <= internal_txelecidle0_ext_pcie;
  --vhdl renameroo for output signals
  txelecidle1_ext_pcie <= internal_txelecidle1_ext_pcie;
  --vhdl renameroo for output signals
  txelecidle2_ext_pcie <= internal_txelecidle2_ext_pcie;
  --vhdl renameroo for output signals
  txelecidle3_ext_pcie <= internal_txelecidle3_ext_pcie;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component pcie_to_hibi_4x_sopc is 
           port (
                 -- 1) global signals:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- the_a2h
                    signal hibi_av_in_to_the_a2h : IN STD_LOGIC;
                    signal hibi_av_out_from_the_a2h : OUT STD_LOGIC;
                    signal hibi_comm_in_to_the_a2h : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal hibi_comm_out_from_the_a2h : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal hibi_data_in_to_the_a2h : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal hibi_data_out_from_the_a2h : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal hibi_empty_in_to_the_a2h : IN STD_LOGIC;
                    signal hibi_full_in_to_the_a2h : IN STD_LOGIC;
                    signal hibi_one_d_in_to_the_a2h : IN STD_LOGIC;
                    signal hibi_one_p_in_to_the_a2h : IN STD_LOGIC;
                    signal hibi_re_out_from_the_a2h : OUT STD_LOGIC;
                    signal hibi_we_out_from_the_a2h : OUT STD_LOGIC;

                 -- the_pcie
                    signal clk125_out_pcie : OUT STD_LOGIC;
                    signal clk250_out_pcie : OUT STD_LOGIC;
                    signal clk500_out_pcie : OUT STD_LOGIC;
                    signal gxb_powerdown_pcie : IN STD_LOGIC;
                    signal pcie_rstn_pcie : IN STD_LOGIC;
                    signal phystatus_ext_pcie : IN STD_LOGIC;
                    signal pipe_mode_pcie : IN STD_LOGIC;
                    signal pll_powerdown_pcie : IN STD_LOGIC;
                    signal powerdown_ext_pcie : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rate_ext_pcie : OUT STD_LOGIC;
                    signal reconfig_clk_pcie : IN STD_LOGIC;
                    signal reconfig_fromgxb_pcie : OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
                    signal reconfig_togxb_pcie : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal refclk_pcie : IN STD_LOGIC;
                    signal rx_in0_pcie : IN STD_LOGIC;
                    signal rx_in1_pcie : IN STD_LOGIC;
                    signal rx_in2_pcie : IN STD_LOGIC;
                    signal rx_in3_pcie : IN STD_LOGIC;
                    signal rxdata0_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata1_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata2_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata3_ext_pcie : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdatak0_ext_pcie : IN STD_LOGIC;
                    signal rxdatak1_ext_pcie : IN STD_LOGIC;
                    signal rxdatak2_ext_pcie : IN STD_LOGIC;
                    signal rxdatak3_ext_pcie : IN STD_LOGIC;
                    signal rxelecidle0_ext_pcie : IN STD_LOGIC;
                    signal rxelecidle1_ext_pcie : IN STD_LOGIC;
                    signal rxelecidle2_ext_pcie : IN STD_LOGIC;
                    signal rxelecidle3_ext_pcie : IN STD_LOGIC;
                    signal rxpolarity0_ext_pcie : OUT STD_LOGIC;
                    signal rxpolarity1_ext_pcie : OUT STD_LOGIC;
                    signal rxpolarity2_ext_pcie : OUT STD_LOGIC;
                    signal rxpolarity3_ext_pcie : OUT STD_LOGIC;
                    signal rxstatus0_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus1_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus2_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus3_ext_pcie : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxvalid0_ext_pcie : IN STD_LOGIC;
                    signal rxvalid1_ext_pcie : IN STD_LOGIC;
                    signal rxvalid2_ext_pcie : IN STD_LOGIC;
                    signal rxvalid3_ext_pcie : IN STD_LOGIC;
                    signal test_in_pcie : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal test_out_pcie : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal tx_out0_pcie : OUT STD_LOGIC;
                    signal tx_out1_pcie : OUT STD_LOGIC;
                    signal tx_out2_pcie : OUT STD_LOGIC;
                    signal tx_out3_pcie : OUT STD_LOGIC;
                    signal txcompl0_ext_pcie : OUT STD_LOGIC;
                    signal txcompl1_ext_pcie : OUT STD_LOGIC;
                    signal txcompl2_ext_pcie : OUT STD_LOGIC;
                    signal txcompl3_ext_pcie : OUT STD_LOGIC;
                    signal txdata0_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata1_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata2_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata3_ext_pcie : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdatak0_ext_pcie : OUT STD_LOGIC;
                    signal txdatak1_ext_pcie : OUT STD_LOGIC;
                    signal txdatak2_ext_pcie : OUT STD_LOGIC;
                    signal txdatak3_ext_pcie : OUT STD_LOGIC;
                    signal txdetectrx_ext_pcie : OUT STD_LOGIC;
                    signal txelecidle0_ext_pcie : OUT STD_LOGIC;
                    signal txelecidle1_ext_pcie : OUT STD_LOGIC;
                    signal txelecidle2_ext_pcie : OUT STD_LOGIC;
                    signal txelecidle3_ext_pcie : OUT STD_LOGIC
                 );
end component pcie_to_hibi_4x_sopc;

component pcie_testbench is 
           port (
                 -- inputs:
                    signal clk125_out : IN STD_LOGIC;
                    signal clk250_out : IN STD_LOGIC;
                    signal clk500_out : IN STD_LOGIC;
                    signal powerdown_ext : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rate_ext : IN STD_LOGIC;
                    signal reconfig_fromgxb : IN STD_LOGIC_VECTOR (16 DOWNTO 0);
                    signal rxpolarity0_ext : IN STD_LOGIC;
                    signal rxpolarity1_ext : IN STD_LOGIC;
                    signal rxpolarity2_ext : IN STD_LOGIC;
                    signal rxpolarity3_ext : IN STD_LOGIC;
                    signal test_out : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal tx_out0 : IN STD_LOGIC;
                    signal tx_out1 : IN STD_LOGIC;
                    signal tx_out2 : IN STD_LOGIC;
                    signal tx_out3 : IN STD_LOGIC;
                    signal txcompl0_ext : IN STD_LOGIC;
                    signal txcompl1_ext : IN STD_LOGIC;
                    signal txcompl2_ext : IN STD_LOGIC;
                    signal txcompl3_ext : IN STD_LOGIC;
                    signal txdata0_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata1_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata2_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdata3_ext : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal txdatak0_ext : IN STD_LOGIC;
                    signal txdatak1_ext : IN STD_LOGIC;
                    signal txdatak2_ext : IN STD_LOGIC;
                    signal txdatak3_ext : IN STD_LOGIC;
                    signal txdetectrx_ext : IN STD_LOGIC;
                    signal txelecidle0_ext : IN STD_LOGIC;
                    signal txelecidle1_ext : IN STD_LOGIC;
                    signal txelecidle2_ext : IN STD_LOGIC;
                    signal txelecidle3_ext : IN STD_LOGIC;

                 -- outputs:
                    signal gxb_powerdown : OUT STD_LOGIC;
                    signal pcie_rstn : OUT STD_LOGIC;
                    signal phystatus_ext : OUT STD_LOGIC;
                    signal pipe_mode : OUT STD_LOGIC;
                    signal pll_powerdown : OUT STD_LOGIC;
                    signal reconfig_clk : OUT STD_LOGIC;
                    signal reconfig_togxb : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal refclk : OUT STD_LOGIC;
                    signal rx_in0 : OUT STD_LOGIC;
                    signal rx_in1 : OUT STD_LOGIC;
                    signal rx_in2 : OUT STD_LOGIC;
                    signal rx_in3 : OUT STD_LOGIC;
                    signal rxdata0_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata1_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata2_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdata3_ext : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rxdatak0_ext : OUT STD_LOGIC;
                    signal rxdatak1_ext : OUT STD_LOGIC;
                    signal rxdatak2_ext : OUT STD_LOGIC;
                    signal rxdatak3_ext : OUT STD_LOGIC;
                    signal rxelecidle0_ext : OUT STD_LOGIC;
                    signal rxelecidle1_ext : OUT STD_LOGIC;
                    signal rxelecidle2_ext : OUT STD_LOGIC;
                    signal rxelecidle3_ext : OUT STD_LOGIC;
                    signal rxstatus0_ext : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus1_ext : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus2_ext : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxstatus3_ext : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal rxvalid0_ext : OUT STD_LOGIC;
                    signal rxvalid1_ext : OUT STD_LOGIC;
                    signal rxvalid2_ext : OUT STD_LOGIC;
                    signal rxvalid3_ext : OUT STD_LOGIC;
                    signal test_in : OUT STD_LOGIC_VECTOR (39 DOWNTO 0)
                 );
end component pcie_testbench;

                signal clk :  STD_LOGIC;
                signal clk125_out_pcie :  STD_LOGIC;
                signal clk250_out_pcie :  STD_LOGIC;
                signal clk500_out_pcie :  STD_LOGIC;
                signal dma_control_port_slave_irq :  STD_LOGIC;
                signal dma_control_port_slave_readyfordata_from_sa :  STD_LOGIC;
                signal dma_read_master_endofpacket :  STD_LOGIC;
                signal dma_write_master_endofpacket :  STD_LOGIC;
                signal gxb_powerdown_pcie :  STD_LOGIC;
                signal hibi_av_in_to_the_a2h :  STD_LOGIC;
                signal hibi_av_out_from_the_a2h :  STD_LOGIC;
                signal hibi_comm_in_to_the_a2h :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal hibi_comm_out_from_the_a2h :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal hibi_data_in_to_the_a2h :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal hibi_data_out_from_the_a2h :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal hibi_empty_in_to_the_a2h :  STD_LOGIC;
                signal hibi_full_in_to_the_a2h :  STD_LOGIC;
                signal hibi_one_d_in_to_the_a2h :  STD_LOGIC;
                signal hibi_one_p_in_to_the_a2h :  STD_LOGIC;
                signal hibi_re_out_from_the_a2h :  STD_LOGIC;
                signal hibi_we_out_from_the_a2h :  STD_LOGIC;
                signal pcie_Control_Register_Access_irq :  STD_LOGIC;
                signal pcie_Rx_Interface_irq :  STD_LOGIC;
                signal pcie_Rx_Interface_irqnumber :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal pcie_rstn_pcie :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_1_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_2_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_3_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcie_to_hibi_4x_sopc_burst_4_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_debugaccess :  STD_LOGIC;
                signal pcie_to_hibi_4x_sopc_burst_5_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal phystatus_ext_pcie :  STD_LOGIC;
                signal pipe_mode_pcie :  STD_LOGIC;
                signal pll_powerdown_pcie :  STD_LOGIC;
                signal powerdown_ext_pcie :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal rate_ext_pcie :  STD_LOGIC;
                signal reconfig_clk_pcie :  STD_LOGIC;
                signal reconfig_fromgxb_pcie :  STD_LOGIC_VECTOR (16 DOWNTO 0);
                signal reconfig_togxb_pcie :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal refclk_pcie :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal rx_in0_pcie :  STD_LOGIC;
                signal rx_in1_pcie :  STD_LOGIC;
                signal rx_in2_pcie :  STD_LOGIC;
                signal rx_in3_pcie :  STD_LOGIC;
                signal rxdata0_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal rxdata1_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal rxdata2_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal rxdata3_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal rxdatak0_ext_pcie :  STD_LOGIC;
                signal rxdatak1_ext_pcie :  STD_LOGIC;
                signal rxdatak2_ext_pcie :  STD_LOGIC;
                signal rxdatak3_ext_pcie :  STD_LOGIC;
                signal rxelecidle0_ext_pcie :  STD_LOGIC;
                signal rxelecidle1_ext_pcie :  STD_LOGIC;
                signal rxelecidle2_ext_pcie :  STD_LOGIC;
                signal rxelecidle3_ext_pcie :  STD_LOGIC;
                signal rxpolarity0_ext_pcie :  STD_LOGIC;
                signal rxpolarity1_ext_pcie :  STD_LOGIC;
                signal rxpolarity2_ext_pcie :  STD_LOGIC;
                signal rxpolarity3_ext_pcie :  STD_LOGIC;
                signal rxstatus0_ext_pcie :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal rxstatus1_ext_pcie :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal rxstatus2_ext_pcie :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal rxstatus3_ext_pcie :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal rxvalid0_ext_pcie :  STD_LOGIC;
                signal rxvalid1_ext_pcie :  STD_LOGIC;
                signal rxvalid2_ext_pcie :  STD_LOGIC;
                signal rxvalid3_ext_pcie :  STD_LOGIC;
                signal test_in_pcie :  STD_LOGIC_VECTOR (39 DOWNTO 0);
                signal test_out_pcie :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal tx_out0_pcie :  STD_LOGIC;
                signal tx_out1_pcie :  STD_LOGIC;
                signal tx_out2_pcie :  STD_LOGIC;
                signal tx_out3_pcie :  STD_LOGIC;
                signal txcompl0_ext_pcie :  STD_LOGIC;
                signal txcompl1_ext_pcie :  STD_LOGIC;
                signal txcompl2_ext_pcie :  STD_LOGIC;
                signal txcompl3_ext_pcie :  STD_LOGIC;
                signal txdata0_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal txdata1_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal txdata2_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal txdata3_ext_pcie :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal txdatak0_ext_pcie :  STD_LOGIC;
                signal txdatak1_ext_pcie :  STD_LOGIC;
                signal txdatak2_ext_pcie :  STD_LOGIC;
                signal txdatak3_ext_pcie :  STD_LOGIC;
                signal txdetectrx_ext_pcie :  STD_LOGIC;
                signal txelecidle0_ext_pcie :  STD_LOGIC;
                signal txelecidle1_ext_pcie :  STD_LOGIC;
                signal txelecidle2_ext_pcie :  STD_LOGIC;
                signal txelecidle3_ext_pcie :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : pcie_to_hibi_4x_sopc
    port map(
      clk125_out_pcie => clk125_out_pcie,
      clk250_out_pcie => clk250_out_pcie,
      clk500_out_pcie => clk500_out_pcie,
      hibi_av_out_from_the_a2h => hibi_av_out_from_the_a2h,
      hibi_comm_out_from_the_a2h => hibi_comm_out_from_the_a2h,
      hibi_data_out_from_the_a2h => hibi_data_out_from_the_a2h,
      hibi_re_out_from_the_a2h => hibi_re_out_from_the_a2h,
      hibi_we_out_from_the_a2h => hibi_we_out_from_the_a2h,
      powerdown_ext_pcie => powerdown_ext_pcie,
      rate_ext_pcie => rate_ext_pcie,
      reconfig_fromgxb_pcie => reconfig_fromgxb_pcie,
      rxpolarity0_ext_pcie => rxpolarity0_ext_pcie,
      rxpolarity1_ext_pcie => rxpolarity1_ext_pcie,
      rxpolarity2_ext_pcie => rxpolarity2_ext_pcie,
      rxpolarity3_ext_pcie => rxpolarity3_ext_pcie,
      test_out_pcie => test_out_pcie,
      tx_out0_pcie => tx_out0_pcie,
      tx_out1_pcie => tx_out1_pcie,
      tx_out2_pcie => tx_out2_pcie,
      tx_out3_pcie => tx_out3_pcie,
      txcompl0_ext_pcie => txcompl0_ext_pcie,
      txcompl1_ext_pcie => txcompl1_ext_pcie,
      txcompl2_ext_pcie => txcompl2_ext_pcie,
      txcompl3_ext_pcie => txcompl3_ext_pcie,
      txdata0_ext_pcie => txdata0_ext_pcie,
      txdata1_ext_pcie => txdata1_ext_pcie,
      txdata2_ext_pcie => txdata2_ext_pcie,
      txdata3_ext_pcie => txdata3_ext_pcie,
      txdatak0_ext_pcie => txdatak0_ext_pcie,
      txdatak1_ext_pcie => txdatak1_ext_pcie,
      txdatak2_ext_pcie => txdatak2_ext_pcie,
      txdatak3_ext_pcie => txdatak3_ext_pcie,
      txdetectrx_ext_pcie => txdetectrx_ext_pcie,
      txelecidle0_ext_pcie => txelecidle0_ext_pcie,
      txelecidle1_ext_pcie => txelecidle1_ext_pcie,
      txelecidle2_ext_pcie => txelecidle2_ext_pcie,
      txelecidle3_ext_pcie => txelecidle3_ext_pcie,
      clk => clk,
      gxb_powerdown_pcie => gxb_powerdown_pcie,
      hibi_av_in_to_the_a2h => hibi_av_in_to_the_a2h,
      hibi_comm_in_to_the_a2h => hibi_comm_in_to_the_a2h,
      hibi_data_in_to_the_a2h => hibi_data_in_to_the_a2h,
      hibi_empty_in_to_the_a2h => hibi_empty_in_to_the_a2h,
      hibi_full_in_to_the_a2h => hibi_full_in_to_the_a2h,
      hibi_one_d_in_to_the_a2h => hibi_one_d_in_to_the_a2h,
      hibi_one_p_in_to_the_a2h => hibi_one_p_in_to_the_a2h,
      pcie_rstn_pcie => pcie_rstn_pcie,
      phystatus_ext_pcie => phystatus_ext_pcie,
      pipe_mode_pcie => pipe_mode_pcie,
      pll_powerdown_pcie => pll_powerdown_pcie,
      reconfig_clk_pcie => reconfig_clk_pcie,
      reconfig_togxb_pcie => reconfig_togxb_pcie,
      refclk_pcie => refclk_pcie,
      reset_n => reset_n,
      rx_in0_pcie => rx_in0_pcie,
      rx_in1_pcie => rx_in1_pcie,
      rx_in2_pcie => rx_in2_pcie,
      rx_in3_pcie => rx_in3_pcie,
      rxdata0_ext_pcie => rxdata0_ext_pcie,
      rxdata1_ext_pcie => rxdata1_ext_pcie,
      rxdata2_ext_pcie => rxdata2_ext_pcie,
      rxdata3_ext_pcie => rxdata3_ext_pcie,
      rxdatak0_ext_pcie => rxdatak0_ext_pcie,
      rxdatak1_ext_pcie => rxdatak1_ext_pcie,
      rxdatak2_ext_pcie => rxdatak2_ext_pcie,
      rxdatak3_ext_pcie => rxdatak3_ext_pcie,
      rxelecidle0_ext_pcie => rxelecidle0_ext_pcie,
      rxelecidle1_ext_pcie => rxelecidle1_ext_pcie,
      rxelecidle2_ext_pcie => rxelecidle2_ext_pcie,
      rxelecidle3_ext_pcie => rxelecidle3_ext_pcie,
      rxstatus0_ext_pcie => rxstatus0_ext_pcie,
      rxstatus1_ext_pcie => rxstatus1_ext_pcie,
      rxstatus2_ext_pcie => rxstatus2_ext_pcie,
      rxstatus3_ext_pcie => rxstatus3_ext_pcie,
      rxvalid0_ext_pcie => rxvalid0_ext_pcie,
      rxvalid1_ext_pcie => rxvalid1_ext_pcie,
      rxvalid2_ext_pcie => rxvalid2_ext_pcie,
      rxvalid3_ext_pcie => rxvalid3_ext_pcie,
      test_in_pcie => test_in_pcie
    );


  --the_pcie_testbench, which is an e_instance
  the_pcie_testbench : pcie_testbench
    port map(
      gxb_powerdown => gxb_powerdown_pcie,
      pcie_rstn => pcie_rstn_pcie,
      phystatus_ext => phystatus_ext_pcie,
      pipe_mode => pipe_mode_pcie,
      pll_powerdown => pll_powerdown_pcie,
      reconfig_clk => reconfig_clk_pcie,
      reconfig_togxb => reconfig_togxb_pcie,
      refclk => refclk_pcie,
      rx_in0 => rx_in0_pcie,
      rx_in1 => rx_in1_pcie,
      rx_in2 => rx_in2_pcie,
      rx_in3 => rx_in3_pcie,
      rxdata0_ext => rxdata0_ext_pcie,
      rxdata1_ext => rxdata1_ext_pcie,
      rxdata2_ext => rxdata2_ext_pcie,
      rxdata3_ext => rxdata3_ext_pcie,
      rxdatak0_ext => rxdatak0_ext_pcie,
      rxdatak1_ext => rxdatak1_ext_pcie,
      rxdatak2_ext => rxdatak2_ext_pcie,
      rxdatak3_ext => rxdatak3_ext_pcie,
      rxelecidle0_ext => rxelecidle0_ext_pcie,
      rxelecidle1_ext => rxelecidle1_ext_pcie,
      rxelecidle2_ext => rxelecidle2_ext_pcie,
      rxelecidle3_ext => rxelecidle3_ext_pcie,
      rxstatus0_ext => rxstatus0_ext_pcie,
      rxstatus1_ext => rxstatus1_ext_pcie,
      rxstatus2_ext => rxstatus2_ext_pcie,
      rxstatus3_ext => rxstatus3_ext_pcie,
      rxvalid0_ext => rxvalid0_ext_pcie,
      rxvalid1_ext => rxvalid1_ext_pcie,
      rxvalid2_ext => rxvalid2_ext_pcie,
      rxvalid3_ext => rxvalid3_ext_pcie,
      test_in => test_in_pcie,
      clk125_out => clk125_out_pcie,
      clk250_out => clk250_out_pcie,
      clk500_out => clk500_out_pcie,
      powerdown_ext => powerdown_ext_pcie,
      rate_ext => rate_ext_pcie,
      reconfig_fromgxb => reconfig_fromgxb_pcie,
      rxpolarity0_ext => rxpolarity0_ext_pcie,
      rxpolarity1_ext => rxpolarity1_ext_pcie,
      rxpolarity2_ext => rxpolarity2_ext_pcie,
      rxpolarity3_ext => rxpolarity3_ext_pcie,
      test_out => test_out_pcie,
      tx_out0 => tx_out0_pcie,
      tx_out1 => tx_out1_pcie,
      tx_out2 => tx_out2_pcie,
      tx_out3 => tx_out3_pcie,
      txcompl0_ext => txcompl0_ext_pcie,
      txcompl1_ext => txcompl1_ext_pcie,
      txcompl2_ext => txcompl2_ext_pcie,
      txcompl3_ext => txcompl3_ext_pcie,
      txdata0_ext => txdata0_ext_pcie,
      txdata1_ext => txdata1_ext_pcie,
      txdata2_ext => txdata2_ext_pcie,
      txdata3_ext => txdata3_ext_pcie,
      txdatak0_ext => txdatak0_ext_pcie,
      txdatak1_ext => txdatak1_ext_pcie,
      txdatak2_ext => txdatak2_ext_pcie,
      txdatak3_ext => txdatak3_ext_pcie,
      txdetectrx_ext => txdetectrx_ext_pcie,
      txelecidle0_ext => txelecidle0_ext_pcie,
      txelecidle1_ext => txelecidle1_ext_pcie,
      txelecidle2_ext => txelecidle2_ext_pcie,
      txelecidle3_ext => txelecidle3_ext_pcie
    );


  process
  begin
    clk <= '0';
    loop
       wait for 5 ns;
       clk <= not clk;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 100 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
