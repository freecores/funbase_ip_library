-- megafunction wizard: %In-System Sources and Probes%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsource_probe 

-- ============================================================
-- File Name: in_sys_sp.vhd
-- Megafunction Name(s):
-- 			altsource_probe
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Build 157 04/27/2011 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;

library altera_mf;
use altera_mf.all;

entity alt_in_sys_sp is
	generic (
	  INSTANCE_INDEX : integer := 0;
    PROBE_WIDTH    : integer := 0;
    SOURCE_WIDTH   : integer := 0 );
  port (
		probe  : in std_logic_vector(PROBE_WIDTH-1 downto 0);
		source : out std_logic_vector(SOURCE_WIDTH-1 downto 0) );
end alt_in_sys_sp;

architecture rtl of alt_in_sys_sp is
  
  component altsource_probe
  generic (
		enable_metastability    : string;
		instance_id             : string;
		probe_width             : natural;
		sld_auto_instance_index : string;
		sld_instance_index      : natural;
		source_initial_value    : string;
		source_width            : natural;
		lpm_type                : string );
	port (
    probe  : in std_logic_vector(PROBE_WIDTH-1 downto 0);
    source : out std_logic_vector(SOURCE_WIDTH-1 downto 0) );
	end component;
  
	signal sub_wire0	: std_logic_vector (0 downto 0);
  
begin
	source    <= sub_wire0(0 downto 0);
  
	altsource_probe_component : altsource_probe
	generic map (
		enable_metastability => "NO",
		instance_id => "NONE",
		probe_width => PROBE_WIDTH,
		sld_auto_instance_index => "YES",
		sld_instance_index => INSTANCE_INDEX,
		source_initial_value => "1",
		source_width => SOURCE_WIDTH,
		lpm_type => "altsource_probe" )
	port map (
		probe => probe,
		source => source );

end rtl;
