-- megafunction wizard: %FIFO%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: dcfifo 

-- ============================================================
-- File Name: fifo_multi_clk.vhd
-- Megafunction Name(s):
-- 			dcfifo
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 10.0 Build 262 08/18/2010 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library altera_mf;
use altera_mf.all;

entity alt_fifo_dc_dw is
	generic ( DATA_WIDTH : integer := 8;
            FIFO_LENGTH : integer := 256;
            CNT_WIDTH : integer := 9;
            
            RDATA_WIDTH : integer := 8;
            RCNT_WIDTH : integer := 9 );
  
  port (
		rclk : in std_logic;
		wclk : in std_logic;
		rst_n : in std_logic;
		
    wdata_in : in std_logic_vector(DATA_WIDTH-1 downto 0);
		rdata_out : out std_logic_vector(RDATA_WIDTH-1 downto 0);
    re_in : in std_logic;
		we_in : in std_logic;
		rempty_out : out std_logic;
		one_d_out : out std_logic;
    two_d_out : out std_logic;
    rcount_out : out std_logic_vector(RCNT_WIDTH-1 downto 0);
		wfull_out : out std_logic;
	  wcount_out : out std_logic_vector(CNT_WIDTH-1 downto 0) );
end alt_fifo_dc_dw;


architecture rtl of alt_fifo_dc_dw is
  
  component dcfifo_mixed_widths
    generic (
    lpm_width               : natural;
    lpm_widthu              : natural;
    lpm_width_r             : natural := 0;
    lpm_widthu_r            : natural := 0;
    lpm_numwords            : natural;
    delay_rdusedw           : natural := 1;
    delay_wrusedw           : natural := 1;
    rdsync_delaypipe        : natural := 0;
    wrsync_delaypipe        : natural := 0;
    intended_device_family  : string := "Stratix";
    lpm_showahead           : string := "OFF";
    underflow_checking      : string := "ON";
    overflow_checking       : string := "ON";
    clocks_are_synchronized : string := "FALSE";
    use_eab                 : string := "ON";
    add_ram_output_register : string := "OFF";
    add_width               : natural := 1;
    ram_block_type          : string := "AUTO";
    add_usedw_msb_bit       : string := "OFF";
    write_aclr_synch        : string := "OFF";
    lpm_hint                : string := "USE_EAB=ON";
    lpm_type                : string := "dcfifo_mixed_widths");
    port (
    data    : in std_logic_vector(lpm_width-1 downto 0);
    rdclk   : in std_logic;
    wrclk   : in std_logic;
    aclr    : in std_logic := '0';
    rdreq   : in std_logic;
    wrreq   : in std_logic;

    rdfull  : out std_logic;
    wrfull  : out std_logic;
    rdempty : out std_logic;
    wrempty : out std_logic;
    rdusedw : out std_logic_vector(lpm_widthu_r-1 downto 0);
    wrusedw : out std_logic_vector(lpm_widthu-1 downto 0);
    q       : out std_logic_vector(lpm_width_r-1 downto 0));
  end component;
  
  signal aclr : std_logic;
  signal rcount : std_logic_vector(RCNT_WIDTH-1 downto 0);

begin
  
  process (rcount)
  begin
    if (rcount = 2) then
      two_d_out <= '1';
      one_d_out <= '0';
    elsif (rcount = 1) then
      one_d_out <= '1';
      two_d_out <= '1';
    else
      one_d_out <= '0';
      two_d_out <= '0';
    end if;
  end process;
  
  aclr <= not(rst_n);
  rcount_out <= rcount;
  
  fifo_0 : dcfifo_mixed_widths
    generic map (
    lpm_width => DATA_WIDTH,
    lpm_widthu => CNT_WIDTH,
    lpm_width_r => RDATA_WIDTH,
    lpm_widthu_r => RCNT_WIDTH,
    lpm_numwords => FIFO_LENGTH,
--    delay_rdusedw => 1,
--    delay_wrusedw => 1,
    rdsync_delaypipe => 4,
    wrsync_delaypipe => 4,
    intended_device_family => "Arria II GX",
    lpm_showahead => "ON",
    underflow_checking => "ON",
    overflow_checking => "ON",
--    clocks_are_synchronized => "FALSE",
    use_eab => "ON",
--    add_ram_output_register => "OFF",
--    add_width => 1,
--    ram_block_type => "AUTO",
    add_usedw_msb_bit => "ON",
    write_aclr_synch => "OFF",
--    lpm_hint => "USE_EAB=ON",
    lpm_type => "dcfifo" )

    port map (
    data => wdata_in,
    rdclk => rclk,
    wrclk => wclk,
    aclr => aclr,
    rdreq => re_in,
    wrreq => we_in,

--    rdfull =>
    wrfull => wfull_out,
    rdempty => rempty_out,
--    wrempty =>
    rdusedw => rcount,
    wrusedw => wcount_out,
    q => rdata_out );
  
end rtl;
