-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt2gxb_reconfig 

-- ============================================================
-- File Name: altpcie_reconfig_3cgx.vhd
-- Megafunction Name(s):
-- 			alt2gxb_reconfig
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 304 01/25/2010 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt2gxb_reconfig CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" ENABLE_BUF_CAL="TRUE" NUMBER_OF_CHANNELS=4 NUMBER_OF_RECONFIG_PORTS=1 RECONFIG_FROMGXB_WIDTH=5 RECONFIG_TOGXB_WIDTH=4 busy reconfig_clk reconfig_fromgxb reconfig_togxb
--VERSION_BEGIN 9.1SP1 cbx_alt2gxb_reconfig 2010:01:25:21:07:46:SJ cbx_alt_cal 2010:01:25:21:07:46:SJ cbx_alt_dprio 2010:01:25:21:07:46:SJ cbx_altsyncram 2010:01:25:21:07:46:SJ cbx_cycloneii 2010:01:25:21:07:46:SJ cbx_lpm_add_sub 2010:01:25:21:07:46:SJ cbx_lpm_compare 2010:01:25:21:07:46:SJ cbx_lpm_counter 2010:01:25:21:07:46:SJ cbx_lpm_decode 2010:01:25:21:07:46:SJ cbx_lpm_mux 2010:01:25:21:07:46:SJ cbx_lpm_shiftreg 2010:01:25:21:07:46:SJ cbx_mgl 2010:01:25:21:15:13:SJ cbx_stratix 2010:01:25:21:07:46:SJ cbx_stratixii 2010:01:25:21:07:46:SJ cbx_stratixiii 2010:01:25:21:07:46:SJ cbx_util_mgl 2010:01:25:21:07:46:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm;

 ARCHITECTURE RTL OF altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm IS

	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  is_adce_all_control :	STD_LOGIC;
	 SIGNAL  is_adce_continuous_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_one_time_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_standby_single_control :	STD_LOGIC;
 BEGIN

	busy <= cal_busy;
	cal_busy <= '0';
	reconfig_togxb <= (OTHERS => '0');

 END RTL; --altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altpcie_reconfig_3cgx IS
	PORT
	(
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		busy		: OUT STD_LOGIC ;
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END altpcie_reconfig_3cgx;


ARCHITECTURE RTL OF altpcie_reconfig_3cgx IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (3 DOWNTO 0);



	COMPONENT altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm
	PORT (
			busy	: OUT STD_LOGIC ;
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	reconfig_togxb    <= sub_wire1(3 DOWNTO 0);

	altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm_component : altpcie_reconfig_3cgx_alt2gxb_reconfig_nlm
	PORT MAP (
		reconfig_clk => reconfig_clk,
		reconfig_fromgxb => reconfig_fromgxb,
		busy => sub_wire0,
		reconfig_togxb => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: PMA NUMERIC "0"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "1"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 INPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 5 0 reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.v TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_inst.v FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_bb.v TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_inst.vhd FALSE
